magic
tech sky130A
magscale 1 2
timestamp 1717184819
<< nwell >>
rect 16843 36653 16901 36672
rect 5462 13550 5580 13580
rect 5462 13490 5648 13550
rect 5462 13464 5580 13490
rect 5460 13444 5586 13464
<< poly >>
rect 4680 14440 4766 14460
rect 4680 14388 4700 14440
rect 4752 14388 4766 14440
rect 4680 14370 4766 14388
rect 6559 14456 6694 14495
rect 6559 14394 6592 14456
rect 6668 14394 6694 14456
rect 4705 14286 4735 14370
rect 6559 14360 6694 14394
rect 6606 14000 6636 14360
rect 6886 12994 6996 13016
rect 6886 12978 6908 12994
rect 6675 12948 6908 12978
rect 6886 12938 6908 12948
rect 6970 12938 6996 12994
rect 6886 12917 6996 12938
rect 6891 12916 6967 12917
rect 4655 11488 4685 12293
rect 4546 11436 4796 11488
rect 4546 11320 4636 11436
rect 4726 11320 4796 11436
rect 4546 11272 4796 11320
<< polycont >>
rect 4700 14388 4752 14440
rect 6592 14394 6668 14456
rect 6908 12938 6970 12994
rect 4636 11320 4726 11436
<< locali >>
rect 16843 36653 16901 36672
rect 4680 14440 4766 14460
rect 4680 14388 4700 14440
rect 4752 14388 4766 14440
rect 4680 14370 4766 14388
rect 6559 14456 6694 14495
rect 6559 14394 6592 14456
rect 6668 14394 6694 14456
rect 6559 14360 6694 14394
rect 5462 13548 5580 13580
rect 5462 13542 5494 13548
rect 5388 13506 5494 13542
rect 5462 13490 5494 13506
rect 5554 13490 5580 13548
rect 5462 13454 5580 13490
rect 6886 12994 6996 13016
rect 6886 12938 6908 12994
rect 6970 12938 6996 12994
rect 3786 12732 3910 12744
rect 3786 12678 3816 12732
rect 3884 12678 3910 12732
rect 3786 12657 3910 12678
rect 4283 12423 4369 12448
rect 4283 12379 4299 12423
rect 4352 12412 4369 12423
rect 4708 12412 4742 12677
rect 4352 12379 4742 12412
rect 4283 12378 4742 12379
rect 4283 12346 4369 12378
rect 5014 11951 5048 12932
rect 6886 12917 6996 12938
rect 6891 12916 6967 12917
rect 4978 11934 5085 11951
rect 4978 11889 5007 11934
rect 5064 11889 5085 11934
rect 4978 11867 5085 11889
rect 1212 11629 1648 11765
rect 1212 11502 1485 11629
rect 1645 11502 1648 11629
rect 5190 11633 5224 12678
rect 5774 11921 5808 12677
rect 5737 11909 5862 11921
rect 5737 11839 5756 11909
rect 5838 11839 5862 11909
rect 5950 11914 5985 12679
rect 6080 12354 6114 12678
rect 6256 12530 6290 12678
rect 6208 12520 6291 12530
rect 6208 12485 6235 12520
rect 6270 12485 6291 12520
rect 6208 12477 6291 12485
rect 6530 12354 6586 12370
rect 6080 12353 6586 12354
rect 6080 12320 6544 12353
rect 6530 12319 6544 12320
rect 6578 12319 6586 12353
rect 6530 12307 6586 12319
rect 5950 11895 6029 11914
rect 5950 11860 5975 11895
rect 6011 11860 6029 11895
rect 5950 11841 6029 11860
rect 5737 11819 5862 11839
rect 5738 11818 5861 11819
rect 5276 11692 5421 11747
rect 5276 11633 5307 11692
rect 5190 11599 5307 11633
rect 5276 11586 5307 11599
rect 5380 11586 5421 11692
rect 5276 11541 5421 11586
rect 4546 11436 4796 11488
rect 4546 11320 4636 11436
rect 4726 11320 4796 11436
rect 4546 11272 4796 11320
rect 1204 10249 1276 10278
rect 1204 10203 1220 10249
rect 1260 10203 1276 10249
rect 1204 10182 1276 10203
rect 1571 5911 1719 5938
rect 1205 5894 1719 5911
rect 1205 5788 1610 5894
rect 1683 5788 1719 5894
rect 1205 5754 1719 5788
rect 1206 4372 1274 5754
rect 1571 5735 1719 5754
rect 11802 4176 11888 4188
rect 11802 4120 11819 4176
rect 11875 4120 11888 4176
rect 11802 4108 11888 4120
rect 1646 3625 2009 3747
rect 1263 3597 2009 3625
rect 1263 3326 1712 3597
rect 1646 3324 1712 3326
rect 1922 3324 2009 3597
rect 1646 3198 2009 3324
rect 10625 1692 11881 1735
rect 10625 1601 10667 1692
rect 10761 1601 11881 1692
rect 10625 1556 11881 1601
<< viali >>
rect 4700 14388 4752 14440
rect 6592 14394 6668 14456
rect 5494 13490 5554 13548
rect 6908 12938 6970 12994
rect 3816 12678 3884 12732
rect 4299 12379 4352 12423
rect 5007 11889 5064 11934
rect 1485 11469 1645 11629
rect 5756 11839 5838 11909
rect 6235 12485 6270 12520
rect 6544 12319 6578 12353
rect 5975 11860 6011 11895
rect 5307 11586 5380 11692
rect 4636 11320 4726 11436
rect 1220 10203 1260 10249
rect 1211 7470 1255 7514
rect 1610 5788 1683 5894
rect 11819 4120 11875 4176
rect 1712 3324 1922 3597
rect 10667 1601 10761 1692
<< metal1 >>
rect 16968 44570 17072 44588
rect 16968 44518 16991 44570
rect 17043 44518 17072 44570
rect 16968 44491 17072 44518
rect 17700 44494 17804 44591
rect 17001 40113 17032 44491
rect 16984 40061 16990 40113
rect 17042 40061 17048 40113
rect 201 38937 501 39037
rect 201 38837 299 38937
rect 399 38934 13817 38937
rect 399 38838 14287 38934
rect 399 38837 13882 38838
rect 201 38737 501 38837
rect 13786 37846 13882 38837
rect 23814 38294 24387 38390
rect 13786 37750 14269 37846
rect 13786 36758 13882 37750
rect 24291 37302 24387 38294
rect 23814 37206 24387 37302
rect 13786 36662 14276 36758
rect 13786 35670 13882 36662
rect 24291 36214 24387 37206
rect 23814 36118 24387 36214
rect 13786 35574 14288 35670
rect 13786 34582 13882 35574
rect 24291 35126 24387 36118
rect 23814 35030 24387 35126
rect 13786 34486 14292 34582
rect 13786 33494 13882 34486
rect 24291 34038 24387 35030
rect 23814 33942 24387 34038
rect 13786 33398 14272 33494
rect 13786 32406 13882 33398
rect 24291 32950 24387 33942
rect 23814 32854 24387 32950
rect 13786 32310 14269 32406
rect 13786 31318 13882 32310
rect 24291 31862 24387 32854
rect 23814 31766 24387 31862
rect 13786 31222 14304 31318
rect 13786 30230 13882 31222
rect 24291 30774 24387 31766
rect 23814 30678 24387 30774
rect 13786 30134 14250 30230
rect 9800 29686 10100 29751
rect 24291 29686 24387 30678
rect 9800 29590 9883 29686
rect 9979 29590 14346 29686
rect 23814 29590 24387 29686
rect 9800 29552 10100 29590
rect 3500 26288 3608 26312
rect 3500 26236 3528 26288
rect 3580 26236 3608 26288
rect 3500 26222 3608 26236
rect 2470 24983 2907 25047
rect 2470 24881 2614 24983
rect 2133 24847 2614 24881
rect 2470 24787 2614 24847
rect 2787 24787 2907 24983
rect 2470 24687 2907 24787
rect 4102 23965 4156 26135
rect 4102 23911 8483 23965
rect 4058 18527 4079 18541
rect 200 16648 500 16682
rect 200 16546 273 16648
rect 411 16625 500 16648
rect 4058 16625 4112 18527
rect 8429 16625 8483 23911
rect 9800 17862 10100 17926
rect 9800 17722 9870 17862
rect 10002 17836 10100 17862
rect 10002 17740 18246 17836
rect 10002 17738 17924 17740
rect 10002 17722 10100 17738
rect 9800 17670 10100 17722
rect 17796 16748 17892 17738
rect 30446 17196 30676 17292
rect 17796 16652 18258 16748
rect 411 16571 8489 16625
rect 411 16570 4099 16571
rect 411 16546 500 16570
rect 200 16505 500 16546
rect 17796 15660 17892 16652
rect 30580 16204 30676 17196
rect 30438 16108 30676 16204
rect 17796 15564 18220 15660
rect 17796 14572 17892 15564
rect 30580 15116 30676 16108
rect 30444 15020 30676 15116
rect 4680 14440 4766 14460
rect 4680 14388 4700 14440
rect 4752 14388 4766 14440
rect 4680 14370 4766 14388
rect 6559 14456 6694 14495
rect 6559 14394 6592 14456
rect 6668 14394 6694 14456
rect 6559 14360 6694 14394
rect 17796 14476 18244 14572
rect 5462 13548 5580 13580
rect 5462 13490 5494 13548
rect 5554 13490 5580 13548
rect 5462 13454 5580 13490
rect 17796 13484 17892 14476
rect 30580 14028 30676 15020
rect 30440 13932 30676 14028
rect 17796 13388 18236 13484
rect 6886 12994 6996 13016
rect 6886 12938 6908 12994
rect 6970 12938 6996 12994
rect 6886 12917 6996 12938
rect 6891 12916 6967 12917
rect 3786 12732 3910 12744
rect 3786 12678 3816 12732
rect 3884 12678 3910 12732
rect 3786 12657 3910 12678
rect 4283 12423 4369 12448
rect 4283 12379 4299 12423
rect 4352 12379 4369 12423
rect 4283 12346 4369 12379
rect 4288 11700 4359 12346
rect 1625 11635 4360 11700
rect 1473 11463 1479 11635
rect 1651 11538 4360 11635
rect 1651 11463 1657 11538
rect 4546 11436 4796 11488
rect 4546 11320 4636 11436
rect 4726 11320 4796 11436
rect 4546 11272 4796 11320
rect 1204 10249 1276 10278
rect 1204 10203 1220 10249
rect 1260 10244 1276 10249
rect 4884 10244 4918 12685
rect 6208 12522 6291 12530
rect 6208 12520 11203 12522
rect 6208 12485 6235 12520
rect 6270 12490 11203 12520
rect 6270 12485 6291 12490
rect 6208 12477 6291 12485
rect 6530 12354 6586 12370
rect 10626 12354 10806 12355
rect 6530 12353 10806 12354
rect 6530 12319 6544 12353
rect 6578 12321 10806 12353
rect 6578 12320 10679 12321
rect 6578 12319 6586 12320
rect 6530 12307 6586 12319
rect 10626 12245 10679 12320
rect 10752 12245 10806 12321
rect 10626 12218 10806 12245
rect 4978 11934 5085 11951
rect 4978 11889 5007 11934
rect 5064 11889 5085 11934
rect 4978 11867 5085 11889
rect 5737 11909 5862 11921
rect 6798 11915 6978 11945
rect 1260 10210 4918 10244
rect 5001 10233 5057 11867
rect 5737 11839 5756 11909
rect 5838 11839 5862 11909
rect 5950 11901 6029 11914
rect 6798 11901 6844 11915
rect 5950 11895 6844 11901
rect 5950 11860 5975 11895
rect 6011 11860 6844 11895
rect 5950 11853 6844 11860
rect 5950 11841 6029 11853
rect 6798 11845 6844 11853
rect 6934 11845 6978 11915
rect 5737 11819 5862 11839
rect 5738 11818 5861 11819
rect 6798 11816 6978 11845
rect 5276 11692 5421 11747
rect 5276 11586 5307 11692
rect 5380 11586 5421 11692
rect 5276 11541 5421 11586
rect 11171 11501 11203 12490
rect 17796 12396 17892 13388
rect 30580 12940 30676 13932
rect 30442 12844 30676 12940
rect 17796 12300 18248 12396
rect 11078 11469 11258 11501
rect 11078 11372 11131 11469
rect 11218 11372 11258 11469
rect 11078 11343 11258 11372
rect 17796 11308 17892 12300
rect 30580 11852 30676 12844
rect 30438 11756 30676 11852
rect 17796 11212 18214 11308
rect 1260 10203 1276 10210
rect 1204 10182 1276 10203
rect 5001 10177 5451 10233
rect 5395 7520 5451 10177
rect 1193 7514 5451 7520
rect 1193 7470 1211 7514
rect 1255 7470 5451 7514
rect 1193 7464 5451 7470
rect 17796 10220 17892 11212
rect 30580 10764 30676 11756
rect 30446 10668 30676 10764
rect 17796 10124 18214 10220
rect 17796 9132 17892 10124
rect 30580 9676 30676 10668
rect 30446 9580 30676 9676
rect 17796 9036 18228 9132
rect 17796 8044 17892 9036
rect 30580 8588 30676 9580
rect 30448 8492 30676 8588
rect 17796 7948 18214 8044
rect 199 7231 501 7258
rect 199 7059 256 7231
rect 444 7183 501 7231
rect 444 7112 11882 7183
rect 444 7059 501 7112
rect 199 7027 501 7059
rect 11811 6884 11882 7112
rect 17796 6956 17892 7948
rect 30580 7500 30676 8492
rect 30438 7404 30676 7500
rect 17796 6860 18430 6956
rect 30580 6930 30676 7404
rect 1571 5894 1719 5938
rect 1571 5788 1610 5894
rect 1683 5788 1719 5894
rect 1571 5735 1719 5788
rect 17796 5868 17892 6860
rect 30580 6834 30868 6930
rect 30772 6412 30868 6834
rect 30434 6316 30868 6412
rect 17796 5772 18236 5868
rect 200 4934 502 5098
rect 200 4762 256 4934
rect 444 4922 502 4934
rect 12243 4922 12339 4923
rect 30772 4922 30868 6316
rect 444 4826 11517 4922
rect 12243 4826 30868 4922
rect 444 4762 502 4826
rect 200 4634 502 4762
rect 11419 4638 11515 4826
rect 12243 4638 12339 4826
rect 11419 4542 12339 4638
rect 11802 4176 11888 4188
rect 11802 4120 11819 4176
rect 11875 4120 11888 4176
rect 11802 4108 11888 4120
rect 1646 3597 2009 3747
rect 1646 3324 1712 3597
rect 1922 3324 2009 3597
rect 1646 3198 2009 3324
rect 10625 1692 10807 1735
rect 10625 1601 10667 1692
rect 10761 1601 10807 1692
rect 10625 1556 10807 1601
rect 16592 1636 16784 1682
rect 16592 1552 16642 1636
rect 16729 1552 16784 1636
rect 16592 1504 16784 1552
<< via1 >>
rect 16991 44518 17043 44570
rect 16990 40061 17042 40113
rect 299 38837 399 38937
rect 9883 29590 9979 29686
rect 3528 26236 3580 26288
rect 2614 24787 2787 24983
rect 273 16546 411 16648
rect 9870 17722 10002 17862
rect 4700 14388 4752 14440
rect 6592 14394 6668 14456
rect 5494 13490 5554 13548
rect 6908 12938 6970 12994
rect 3816 12678 3884 12732
rect 1479 11629 1651 11635
rect 1479 11469 1485 11629
rect 1485 11469 1645 11629
rect 1645 11469 1651 11629
rect 1479 11463 1651 11469
rect 4636 11320 4726 11436
rect 10679 12245 10752 12321
rect 5756 11839 5838 11909
rect 6844 11845 6934 11915
rect 5307 11586 5380 11692
rect 11131 11372 11218 11469
rect 256 7059 444 7231
rect 1610 5788 1683 5894
rect 256 4762 444 4934
rect 11819 4120 11875 4176
rect 1712 3324 1922 3597
rect 10667 1601 10761 1692
rect 16642 1552 16729 1636
<< metal2 >>
rect 16987 44574 17047 44583
rect 17721 44575 17781 44584
rect 16985 44518 16987 44570
rect 17047 44518 17049 44570
rect 16987 44505 17047 44514
rect 17721 44506 17781 44515
rect 991 42341 1135 42354
rect 991 42285 1028 42341
rect 1091 42325 1135 42341
rect 17723 42325 17779 44506
rect 31442 44285 31571 44291
rect 29461 44165 29470 44285
rect 29590 44280 31571 44285
rect 29590 44170 31450 44280
rect 31560 44170 31571 44280
rect 29590 44165 31571 44170
rect 31442 44160 31571 44165
rect 28721 43912 28865 43924
rect 31193 43912 31323 43918
rect 28721 43792 28732 43912
rect 28852 43907 31323 43912
rect 28852 43797 31201 43907
rect 31311 43797 31323 43907
rect 28852 43792 31323 43797
rect 28721 43781 28865 43792
rect 31193 43787 31323 43792
rect 27984 43476 28128 43488
rect 30721 43476 30851 43481
rect 27984 43356 27996 43476
rect 28116 43471 30851 43476
rect 28116 43361 30730 43471
rect 30840 43361 30851 43471
rect 28116 43356 30851 43361
rect 27984 43345 28128 43356
rect 30721 43350 30851 43356
rect 27253 43143 27397 43154
rect 30768 43143 30898 43149
rect 27253 43023 27264 43143
rect 27384 43138 30898 43143
rect 27384 43028 30778 43138
rect 30888 43028 30898 43138
rect 27384 43023 30898 43028
rect 27253 43011 27397 43023
rect 30768 43018 30898 43023
rect 1091 42285 22144 42325
rect 991 42269 22144 42285
rect 991 42266 1135 42269
rect 695 41555 809 41565
rect 695 41498 723 41555
rect 782 41553 809 41555
rect 782 41498 16164 41553
rect 22088 41503 22144 42269
rect 695 41497 16164 41498
rect 695 41481 809 41497
rect 16990 40113 17042 40119
rect 16120 40071 16990 40102
rect 16990 40055 17042 40061
rect 201 38937 501 39037
rect 201 38837 299 38937
rect 399 38837 501 38937
rect 201 38737 501 38837
rect 9800 29686 10100 29751
rect 9800 29590 9883 29686
rect 9979 29590 10100 29686
rect 9800 29552 10100 29590
rect 16039 27989 16252 28007
rect 16039 27819 16060 27989
rect 16230 27819 16252 27989
rect 16039 27790 16252 27819
rect 22036 27964 22216 27990
rect 22036 27852 22075 27964
rect 22177 27852 22216 27964
rect 22036 27810 22216 27852
rect 17626 27175 30412 27180
rect 17622 27065 17631 27175
rect 17741 27065 30412 27175
rect 17626 27060 30412 27065
rect 30532 27060 30541 27180
rect 3500 26288 3608 26312
rect 3500 26236 3528 26288
rect 3580 26236 3608 26288
rect 3500 26222 3608 26236
rect 2470 24983 2907 25047
rect 2470 24787 2614 24983
rect 2787 24787 2907 24983
rect 2470 24687 2907 24787
rect 3524 24231 3582 26222
rect 9263 24442 9424 24485
rect 9263 24382 9313 24442
rect 9373 24382 9424 24442
rect 9263 24325 9424 24382
rect 9314 24231 9372 24325
rect 3524 24173 20783 24231
rect 20725 21864 20783 24173
rect 20698 21858 20808 21864
rect 20698 21802 20728 21858
rect 20786 21802 20808 21858
rect 20698 21780 20808 21802
rect 14492 21442 27946 21494
rect 3882 17014 3934 18624
rect 8862 17854 9023 17903
rect 8862 17794 8917 17854
rect 8977 17794 9023 17854
rect 8862 17743 9023 17794
rect 9800 17862 10100 17926
rect 8921 17014 8973 17743
rect 9800 17722 9870 17862
rect 10002 17722 10100 17862
rect 9800 17670 10100 17722
rect 14492 17014 14544 21442
rect 3882 16962 14544 17014
rect 17626 20483 17746 20492
rect 20654 20458 20838 20492
rect 20654 20396 20708 20458
rect 20778 20396 20838 20458
rect 20654 20370 20838 20396
rect 200 16648 500 16682
rect 200 16546 273 16648
rect 411 16546 500 16648
rect 200 16505 500 16546
rect 2916 14490 4754 14542
rect 200 12796 500 12824
rect 200 12738 1650 12796
rect 200 12580 264 12738
rect 388 12580 1650 12738
rect 200 12540 1650 12580
rect 200 12520 500 12540
rect 1479 11635 1651 11641
rect 1479 11457 1651 11463
rect 2916 9878 2968 14490
rect 4702 14460 4754 14490
rect 4680 14440 4766 14460
rect 4680 14388 4700 14440
rect 4752 14388 4766 14440
rect 4680 14370 4766 14388
rect 6559 14456 6694 14495
rect 6559 14394 6592 14456
rect 6668 14394 6694 14456
rect 6559 14360 6694 14394
rect 9798 13954 10102 14044
rect 8526 13936 10102 13954
rect 8526 13778 9894 13936
rect 10018 13778 10102 13936
rect 8526 13730 10102 13778
rect 9798 13688 10102 13730
rect 5462 13548 5580 13580
rect 5462 13490 5494 13548
rect 5554 13490 5580 13548
rect 5462 13454 5580 13490
rect 6886 12994 6996 13016
rect 6886 12938 6908 12994
rect 6970 12938 6996 12994
rect 6886 12917 6996 12938
rect 6891 12916 6967 12917
rect 3786 12732 3910 12744
rect 3786 12678 3816 12732
rect 3884 12678 3910 12732
rect 3786 12657 3910 12678
rect 10626 12321 10806 12355
rect 10626 12245 10679 12321
rect 10752 12245 10806 12321
rect 10626 12219 10806 12245
rect 5737 11909 5862 11921
rect 5737 11839 5756 11909
rect 5838 11839 5862 11909
rect 5737 11819 5862 11839
rect 6798 11915 6978 11945
rect 6798 11845 6844 11915
rect 6934 11845 6978 11915
rect 5738 11818 5861 11819
rect 6798 11816 6978 11845
rect 5276 11692 5429 11747
rect 5276 11586 5307 11692
rect 5380 11687 5429 11692
rect 5380 11608 5933 11687
rect 5380 11586 5429 11608
rect 5276 11541 5429 11586
rect 4546 11436 4796 11488
rect 4546 11320 4636 11436
rect 4726 11320 4796 11436
rect 4546 11272 4796 11320
rect 4612 10034 5152 10100
rect 4612 9878 4726 10034
rect 2916 9826 4726 9878
rect 4612 9786 4726 9826
rect 5044 9786 5152 10034
rect 4612 9712 5152 9786
rect 199 7231 501 7258
rect 199 7059 256 7231
rect 444 7059 501 7231
rect 199 7027 501 7059
rect 1571 5916 1719 5938
rect 5795 5916 5933 11608
rect 11078 11469 11258 11501
rect 11078 11372 11131 11469
rect 11218 11372 11258 11469
rect 11078 11343 11258 11372
rect 17626 7858 17746 20363
rect 20714 20180 20770 20370
rect 27890 20230 27946 21442
rect 17621 7847 17758 7858
rect 17621 7737 17631 7847
rect 17741 7737 17758 7847
rect 17621 7725 17758 7737
rect 1571 5894 5933 5916
rect 1571 5788 1610 5894
rect 1683 5788 5933 5894
rect 1571 5778 5933 5788
rect 1571 5735 1719 5778
rect 200 4934 502 5098
rect 200 4762 256 4934
rect 444 4762 502 4934
rect 200 4634 502 4762
rect 11802 4176 11888 4188
rect 11802 4120 11819 4176
rect 11875 4120 11888 4176
rect 11802 4108 11888 4120
rect 1646 3597 2009 3747
rect 1646 3324 1712 3597
rect 1922 3324 2009 3597
rect 1646 3198 2009 3324
rect 14230 3133 14391 3203
rect 14230 3073 14269 3133
rect 14329 3131 14391 3133
rect 18046 3131 18102 3700
rect 14329 3075 18102 3131
rect 14329 3073 14391 3075
rect 14230 3043 14391 3073
rect 13954 2992 14058 3009
rect 13954 2932 13977 2992
rect 14037 2990 14058 2992
rect 19610 2990 19666 3728
rect 14037 2934 19666 2990
rect 14037 2932 14058 2934
rect 13954 2912 14058 2932
rect 13715 2810 13819 2830
rect 13715 2750 13736 2810
rect 13796 2808 13819 2810
rect 21174 2808 21230 3714
rect 13796 2752 21230 2808
rect 13796 2750 13819 2752
rect 13715 2733 13819 2750
rect 13522 2678 13626 2696
rect 13522 2618 13545 2678
rect 13605 2676 13626 2678
rect 22738 2676 22794 3728
rect 13605 2620 22794 2676
rect 13605 2618 13626 2620
rect 13522 2599 13626 2618
rect 13331 2560 13435 2577
rect 13331 2500 13354 2560
rect 13414 2558 13435 2560
rect 24302 2558 24358 3705
rect 13414 2502 24358 2558
rect 13414 2500 13435 2502
rect 13331 2480 13435 2500
rect 13125 2400 13229 2420
rect 13125 2340 13149 2400
rect 13209 2398 13229 2400
rect 25866 2398 25922 3700
rect 13209 2342 25922 2398
rect 13209 2340 13229 2342
rect 13125 2323 13229 2340
rect 12930 2251 13034 2267
rect 12930 2191 12952 2251
rect 13012 2249 13034 2251
rect 27430 2249 27486 3775
rect 13012 2193 27486 2249
rect 13012 2191 13034 2193
rect 12930 2170 13034 2191
rect 12728 2036 12832 2054
rect 12728 1976 12752 2036
rect 12812 2034 12832 2036
rect 28994 2034 29050 3751
rect 12812 1978 29050 2034
rect 12812 1976 12832 1978
rect 12728 1957 12832 1976
rect 12488 1882 12592 1900
rect 12488 1822 12508 1882
rect 12568 1880 12592 1882
rect 30558 1880 30614 3740
rect 12568 1824 30614 1880
rect 12568 1822 12592 1824
rect 12488 1803 12592 1822
rect 10625 1692 10807 1735
rect 10625 1601 10667 1692
rect 10761 1601 10807 1692
rect 16592 1636 16784 1682
rect 16592 1628 16642 1636
rect 10625 1556 10807 1601
rect 12392 1567 16642 1628
rect 4785 1454 4966 1496
rect 4785 1383 4836 1454
rect 4910 1408 4966 1454
rect 12392 1408 12453 1567
rect 16592 1552 16642 1567
rect 16729 1552 16784 1636
rect 16592 1504 16784 1552
rect 4910 1383 12453 1408
rect 4785 1348 12453 1383
rect 4791 1347 12453 1348
<< via2 >>
rect 16987 44570 17047 44574
rect 16987 44518 16991 44570
rect 16991 44518 17043 44570
rect 17043 44518 17047 44570
rect 16987 44514 17047 44518
rect 17721 44515 17781 44575
rect 1028 42285 1091 42341
rect 29470 44165 29590 44285
rect 31450 44170 31560 44280
rect 28732 43792 28852 43912
rect 31201 43797 31311 43907
rect 27996 43356 28116 43476
rect 30730 43361 30840 43471
rect 27264 43023 27384 43143
rect 30778 43028 30888 43138
rect 723 41498 782 41555
rect 299 38837 399 38937
rect 9883 29590 9979 29686
rect 16060 27819 16230 27989
rect 22075 27852 22177 27964
rect 17631 27065 17741 27175
rect 30412 27060 30532 27180
rect 2614 24787 2787 24983
rect 9313 24382 9373 24442
rect 20728 21802 20786 21858
rect 8917 17794 8977 17854
rect 9870 17722 10002 17862
rect 17626 20363 17746 20483
rect 20708 20396 20778 20458
rect 273 16546 411 16648
rect 264 12580 388 12738
rect 6592 14394 6668 14456
rect 9894 13778 10018 13936
rect 5494 13490 5554 13548
rect 6908 12938 6970 12994
rect 10679 12245 10752 12321
rect 5756 11839 5838 11909
rect 6844 11845 6934 11915
rect 4636 11320 4726 11436
rect 4726 9786 5044 10034
rect 256 7059 444 7231
rect 11131 11372 11218 11469
rect 17631 7737 17741 7847
rect 256 4762 444 4934
rect 11819 4120 11875 4176
rect 1712 3324 1922 3597
rect 14269 3073 14329 3133
rect 13977 2932 14037 2992
rect 13736 2750 13796 2810
rect 13545 2618 13605 2678
rect 13354 2500 13414 2560
rect 13149 2340 13209 2400
rect 12952 2191 13012 2251
rect 12752 1976 12812 2036
rect 12508 1822 12568 1882
rect 10667 1601 10761 1692
rect 4836 1383 4910 1454
rect 16642 1552 16729 1636
<< metal3 >>
rect 30856 44763 31216 44809
rect 30856 44626 30956 44763
rect 31070 44626 31216 44763
rect 16968 44579 17072 44588
rect 16968 44509 16982 44579
rect 17052 44509 17072 44579
rect 16968 44491 17072 44509
rect 17700 44580 17804 44591
rect 17700 44510 17716 44580
rect 17786 44510 17804 44580
rect 30856 44549 31216 44626
rect 17700 44494 17804 44510
rect 29465 44290 29595 44296
rect 14041 44171 14105 44177
rect 13313 44163 13377 44169
rect 29465 44165 29470 44170
rect 29590 44165 29595 44170
rect 29465 44160 29595 44165
rect 14041 44101 14105 44107
rect 13313 44093 13377 44099
rect 9305 43781 9311 43845
rect 9375 43843 9381 43845
rect 13315 43843 13375 44093
rect 9375 43783 13375 43843
rect 9375 43781 9381 43783
rect 8909 43523 8915 43587
rect 8979 43585 8985 43587
rect 14043 43585 14103 44101
rect 28721 43917 28865 43924
rect 28721 43787 28727 43917
rect 28857 43787 28865 43917
rect 28721 43781 28865 43787
rect 8979 43525 14103 43585
rect 8979 43523 8985 43525
rect 27984 43481 28128 43488
rect 27984 43351 27991 43481
rect 28121 43351 28128 43481
rect 27984 43345 28128 43351
rect 30721 43475 30851 43481
rect 30721 43357 30726 43475
rect 30844 43357 30851 43475
rect 30721 43350 30851 43357
rect 27253 43148 27397 43154
rect 27253 43018 27259 43148
rect 27389 43018 27397 43148
rect 30768 43142 30898 43149
rect 30768 43024 30774 43142
rect 30892 43024 30898 43142
rect 30768 43018 30898 43024
rect 27253 43011 27397 43018
rect 821 42726 910 42733
rect 821 42659 840 42726
rect 904 42721 910 42726
rect 12555 42728 12671 42734
rect 12555 42721 12581 42728
rect 904 42664 12581 42721
rect 12645 42664 12671 42728
rect 904 42659 12671 42664
rect 821 42658 12671 42659
rect 821 42653 910 42658
rect 12555 42647 12671 42658
rect 991 42341 1135 42354
rect 991 42285 1028 42341
rect 1091 42285 1135 42341
rect 991 42266 1135 42285
rect 695 41555 809 41565
rect 695 41498 723 41555
rect 782 41498 809 41555
rect 695 41481 809 41498
rect 201 38942 501 39037
rect 201 38832 294 38942
rect 404 38832 501 38942
rect 201 38737 501 38832
rect 200 16648 500 16682
rect 200 16546 273 16648
rect 411 16546 500 16648
rect 200 16505 500 16546
rect 713 13221 774 41481
rect 1011 14715 1085 42266
rect 30964 42055 31085 44549
rect 31445 44284 31565 44285
rect 31440 44166 31446 44284
rect 31564 44166 31570 44284
rect 31445 44165 31565 44166
rect 31193 43911 31323 43918
rect 31191 43793 31197 43911
rect 31315 43793 31323 43911
rect 31193 43787 31323 43793
rect 10923 41934 31085 42055
rect 2840 31963 8299 32159
rect 2840 25047 3036 31963
rect 2470 24983 3036 25047
rect 2470 24787 2614 24983
rect 2787 24788 3036 24983
rect 8103 25086 8299 31963
rect 10923 30855 11044 41934
rect 13459 37807 13465 37871
rect 13529 37869 13535 37871
rect 13529 37809 13615 37869
rect 13529 37807 13535 37809
rect 24952 37806 25789 37926
rect 25909 37806 25915 37926
rect 10923 30734 13261 30855
rect 24961 30734 26508 30854
rect 26628 30734 26634 30854
rect 9800 29691 10100 29751
rect 9800 29585 9878 29691
rect 9984 29585 10100 29691
rect 9800 29552 10100 29585
rect 12998 25702 13118 30734
rect 16039 27993 16252 28007
rect 16039 27815 16056 27993
rect 16234 27815 16252 27993
rect 16039 27790 16252 27815
rect 22036 27964 22216 27990
rect 22036 27852 22075 27964
rect 22177 27852 22216 27964
rect 22036 27810 22216 27852
rect 30407 27180 30537 27185
rect 17626 27175 17746 27180
rect 17626 27065 17631 27175
rect 17741 27065 17746 27175
rect 12998 25582 16710 25702
rect 15718 25086 16086 25137
rect 8103 25063 16086 25086
rect 8103 24901 15803 25063
rect 15995 24901 16086 25063
rect 8103 24890 16086 24901
rect 15718 24810 16086 24890
rect 2787 24787 2907 24788
rect 2470 24687 2907 24787
rect 9263 24447 9424 24485
rect 9263 24377 9308 24447
rect 9378 24377 9424 24447
rect 9263 24325 9424 24377
rect 8862 17859 9023 17903
rect 8862 17789 8912 17859
rect 8982 17789 9023 17859
rect 8862 17743 9023 17789
rect 9800 17862 10100 17926
rect 9800 17722 9870 17862
rect 10002 17722 10100 17862
rect 9800 17670 10100 17722
rect 16590 16012 16710 25582
rect 17626 20488 17746 27065
rect 30407 27175 30412 27180
rect 30532 27175 30537 27180
rect 30407 27049 30537 27055
rect 20698 21858 20808 21864
rect 20698 21802 20728 21858
rect 20786 21802 20808 21858
rect 20698 21780 20808 21802
rect 20724 20492 20794 21780
rect 17621 20483 17751 20488
rect 17621 20363 17626 20483
rect 17746 20363 17751 20483
rect 20654 20458 20838 20492
rect 20654 20396 20708 20458
rect 20778 20396 20838 20458
rect 20654 20370 20838 20396
rect 17621 20358 17751 20363
rect 16590 15892 17252 16012
rect 1011 14641 6666 14715
rect 6592 14530 6666 14641
rect 6592 14495 6668 14530
rect 6559 14456 6694 14495
rect 6559 14394 6592 14456
rect 6668 14394 6694 14456
rect 6559 14360 6694 14394
rect 9798 13936 10102 14044
rect 9798 13778 9894 13936
rect 10018 13778 10102 13936
rect 9798 13688 10102 13778
rect 30982 13836 31102 13842
rect 30982 13710 31102 13716
rect 5462 13550 5580 13580
rect 5462 13548 6458 13550
rect 5462 13490 5494 13548
rect 5554 13490 6458 13548
rect 5462 13454 5580 13490
rect 6398 13221 6458 13490
rect 713 13160 6970 13221
rect 200 12738 500 12824
rect 200 12580 264 12738
rect 388 12580 500 12738
rect 200 12520 500 12580
rect 5737 11909 5862 11921
rect 5737 11839 5756 11909
rect 5838 11839 5862 11909
rect 5737 11819 5862 11839
rect 5738 11818 5861 11819
rect 4612 10034 5152 10100
rect 4612 9786 4726 10034
rect 5044 9786 5152 10034
rect 4612 9712 5152 9786
rect 199 7231 501 7258
rect 199 7059 256 7231
rect 444 7059 501 7231
rect 199 7027 501 7059
rect 200 4934 502 5098
rect 200 4762 256 4934
rect 444 4762 502 4934
rect 200 4634 502 4762
rect 6398 4177 6458 13160
rect 6909 13055 6970 13160
rect 6908 13016 6970 13055
rect 6886 12994 6996 13016
rect 6886 12938 6908 12994
rect 6970 12938 6996 12994
rect 6886 12917 6996 12938
rect 6891 12916 6967 12917
rect 10626 12321 10806 12355
rect 10626 12245 10679 12321
rect 10752 12245 10806 12321
rect 10626 12219 10806 12245
rect 6798 11915 6978 11945
rect 6798 11845 6844 11915
rect 6934 11845 6978 11915
rect 6798 11816 6978 11845
rect 11078 11469 11258 11501
rect 11078 11372 11131 11469
rect 11218 11372 11258 11469
rect 11078 11343 11258 11372
rect 17626 7847 17746 7852
rect 17626 7737 17631 7847
rect 17741 7737 17746 7847
rect 17626 7732 17746 7737
rect 31440 5676 31571 5683
rect 31440 5556 31445 5676
rect 31565 5556 31571 5676
rect 31440 5550 31571 5556
rect 11802 4177 11888 4188
rect 6398 4176 11888 4177
rect 6398 4120 11819 4176
rect 11875 4120 11888 4176
rect 6398 4117 11888 4120
rect 11802 4108 11888 4117
rect 1646 3613 2009 3747
rect 9800 3613 10099 3614
rect 1646 3597 10099 3613
rect 1646 3324 1712 3597
rect 1922 3546 10099 3597
rect 1922 3363 9875 3546
rect 10044 3363 10099 3546
rect 1922 3324 10099 3363
rect 1646 3315 10099 3324
rect 1646 3314 10046 3315
rect 1646 3198 2009 3314
rect 14230 3138 14391 3203
rect 14230 3068 14264 3138
rect 14334 3068 14391 3138
rect 14230 3043 14391 3068
rect 13954 2997 14058 3009
rect 13954 2927 13972 2997
rect 14042 2927 14058 2997
rect 13954 2912 14058 2927
rect 13715 2815 13819 2830
rect 13715 2745 13731 2815
rect 13801 2745 13819 2815
rect 13715 2733 13819 2745
rect 13522 2683 13626 2696
rect 13522 2613 13540 2683
rect 13610 2613 13626 2683
rect 13522 2599 13626 2613
rect 13331 2565 13435 2577
rect 13331 2495 13349 2565
rect 13419 2495 13435 2565
rect 13331 2480 13435 2495
rect 13125 2405 13229 2420
rect 13125 2335 13144 2405
rect 13214 2335 13229 2405
rect 13125 2323 13229 2335
rect 12930 2256 13034 2267
rect 12930 2186 12947 2256
rect 13017 2186 13034 2256
rect 12930 2170 13034 2186
rect 12728 2041 12832 2054
rect 12728 1971 12747 2041
rect 12817 1971 12832 2041
rect 12728 1957 12832 1971
rect 12488 1887 12592 1900
rect 12488 1817 12503 1887
rect 12573 1817 12592 1887
rect 12488 1803 12592 1817
rect 10625 1692 10807 1735
rect 10625 1601 10667 1692
rect 10761 1601 10807 1692
rect 10625 1556 10807 1601
rect 16589 1636 16786 1685
rect 16589 1552 16642 1636
rect 16729 1552 16786 1636
rect 16589 1504 16786 1552
rect 4785 1454 4967 1496
rect 4785 1383 4836 1454
rect 4910 1383 4967 1454
rect 4785 1346 4967 1383
rect 16188 1247 16424 1296
rect 2674 1243 16424 1247
rect 2674 1242 16248 1243
rect 2674 1177 2737 1242
rect 2801 1177 16248 1242
rect 2674 1155 16248 1177
rect 16188 1151 16248 1155
rect 16346 1151 16424 1243
rect 16188 1115 16424 1151
<< rmetal3 >>
rect 4546 11436 4796 11488
rect 4546 11320 4636 11436
rect 4726 11320 4796 11436
rect 4546 11272 4796 11320
<< via3 >>
rect 30956 44626 31070 44763
rect 16982 44574 17052 44579
rect 16982 44514 16987 44574
rect 16987 44514 17047 44574
rect 17047 44514 17052 44574
rect 16982 44509 17052 44514
rect 17716 44575 17786 44580
rect 17716 44515 17721 44575
rect 17721 44515 17781 44575
rect 17781 44515 17786 44575
rect 17716 44510 17786 44515
rect 29465 44285 29595 44290
rect 13313 44099 13377 44163
rect 14041 44107 14105 44171
rect 29465 44170 29470 44285
rect 29470 44170 29590 44285
rect 29590 44170 29595 44285
rect 9311 43781 9375 43845
rect 8915 43523 8979 43587
rect 28727 43912 28857 43917
rect 28727 43792 28732 43912
rect 28732 43792 28852 43912
rect 28852 43792 28857 43912
rect 28727 43787 28857 43792
rect 27991 43476 28121 43481
rect 27991 43356 27996 43476
rect 27996 43356 28116 43476
rect 28116 43356 28121 43476
rect 27991 43351 28121 43356
rect 30726 43471 30844 43475
rect 30726 43361 30730 43471
rect 30730 43361 30840 43471
rect 30840 43361 30844 43471
rect 30726 43357 30844 43361
rect 27259 43143 27389 43148
rect 27259 43023 27264 43143
rect 27264 43023 27384 43143
rect 27384 43023 27389 43143
rect 27259 43018 27389 43023
rect 30774 43138 30892 43142
rect 30774 43028 30778 43138
rect 30778 43028 30888 43138
rect 30888 43028 30892 43138
rect 30774 43024 30892 43028
rect 840 42659 904 42726
rect 12581 42664 12645 42728
rect 294 38937 404 38942
rect 294 38837 299 38937
rect 299 38837 399 38937
rect 399 38837 404 38937
rect 294 38832 404 38837
rect 273 16546 411 16648
rect 31446 44280 31564 44284
rect 31446 44170 31450 44280
rect 31450 44170 31560 44280
rect 31560 44170 31564 44280
rect 31446 44166 31564 44170
rect 31197 43907 31315 43911
rect 31197 43797 31201 43907
rect 31201 43797 31311 43907
rect 31311 43797 31315 43907
rect 31197 43793 31315 43797
rect 13465 37807 13529 37871
rect 25789 37806 25909 37926
rect 26508 30734 26628 30854
rect 9878 29686 9984 29691
rect 9878 29590 9883 29686
rect 9883 29590 9979 29686
rect 9979 29590 9984 29686
rect 9878 29585 9984 29590
rect 16056 27989 16234 27993
rect 16056 27819 16060 27989
rect 16060 27819 16230 27989
rect 16230 27819 16234 27989
rect 16056 27815 16234 27819
rect 22075 27852 22177 27964
rect 15803 24901 15995 25063
rect 9308 24442 9378 24447
rect 9308 24382 9313 24442
rect 9313 24382 9373 24442
rect 9373 24382 9378 24442
rect 9308 24377 9378 24382
rect 8912 17854 8982 17859
rect 8912 17794 8917 17854
rect 8917 17794 8977 17854
rect 8977 17794 8982 17854
rect 8912 17789 8982 17794
rect 9870 17722 10002 17862
rect 30407 27060 30412 27175
rect 30412 27060 30532 27175
rect 30532 27060 30537 27175
rect 30407 27055 30537 27060
rect 30773 17796 30893 17916
rect 9894 13778 10018 13936
rect 30982 13716 31102 13836
rect 264 12580 388 12738
rect 5756 11839 5838 11909
rect 4636 11320 4726 11436
rect 4726 9786 5044 10034
rect 256 7059 444 7231
rect 256 4762 444 4934
rect 10679 12245 10752 12321
rect 6844 11845 6934 11915
rect 11131 11372 11218 11469
rect 31196 9636 31316 9756
rect 31445 5556 31565 5676
rect 9875 3363 10044 3546
rect 14264 3133 14334 3138
rect 14264 3073 14269 3133
rect 14269 3073 14329 3133
rect 14329 3073 14334 3133
rect 14264 3068 14334 3073
rect 13972 2992 14042 2997
rect 13972 2932 13977 2992
rect 13977 2932 14037 2992
rect 14037 2932 14042 2992
rect 13972 2927 14042 2932
rect 13731 2810 13801 2815
rect 13731 2750 13736 2810
rect 13736 2750 13796 2810
rect 13796 2750 13801 2810
rect 13731 2745 13801 2750
rect 13540 2678 13610 2683
rect 13540 2618 13545 2678
rect 13545 2618 13605 2678
rect 13605 2618 13610 2678
rect 13540 2613 13610 2618
rect 13349 2560 13419 2565
rect 13349 2500 13354 2560
rect 13354 2500 13414 2560
rect 13414 2500 13419 2560
rect 13349 2495 13419 2500
rect 13144 2400 13214 2405
rect 13144 2340 13149 2400
rect 13149 2340 13209 2400
rect 13209 2340 13214 2400
rect 13144 2335 13214 2340
rect 12947 2251 13017 2256
rect 12947 2191 12952 2251
rect 12952 2191 13012 2251
rect 13012 2191 13017 2251
rect 12947 2186 13017 2191
rect 12747 2036 12817 2041
rect 12747 1976 12752 2036
rect 12752 1976 12812 2036
rect 12812 1976 12817 2036
rect 12747 1971 12817 1976
rect 12503 1882 12573 1887
rect 12503 1822 12508 1882
rect 12508 1822 12568 1882
rect 12568 1822 12573 1882
rect 12503 1817 12573 1822
rect 10667 1601 10761 1692
rect 16642 1552 16729 1636
rect 4836 1383 4910 1454
rect 2737 1177 2801 1242
rect 16248 1151 16346 1243
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44888 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 200 39037 500 44152
rect 9310 43845 9376 43846
rect 9310 43781 9311 43845
rect 9375 43781 9376 43845
rect 9310 43780 9376 43781
rect 8914 43587 8980 43588
rect 8914 43523 8915 43587
rect 8979 43523 8980 43587
rect 8914 43522 8980 43523
rect 821 42726 910 42733
rect 821 42659 840 42726
rect 904 42659 910 42726
rect 821 42653 910 42659
rect 200 38942 501 39037
rect 200 38832 294 38942
rect 404 38832 501 38942
rect 200 38737 501 38832
rect 200 16648 500 38737
rect 200 16546 273 16648
rect 411 16546 500 16648
rect 200 12738 500 16546
rect 200 12580 264 12738
rect 388 12580 500 12738
rect 200 7258 500 12580
rect 842 11893 904 42653
rect 8917 17903 8977 43522
rect 9313 24485 9373 43780
rect 9800 29691 10100 44152
rect 12574 42734 12634 45152
rect 13310 45010 13370 45152
rect 13310 44952 13375 45010
rect 14046 44978 14106 45152
rect 13315 44164 13375 44952
rect 14043 44952 14106 44978
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44980 17050 45152
rect 17726 45026 17786 45152
rect 16987 44952 17050 44980
rect 17721 44952 17786 45026
rect 18462 45006 18522 45152
rect 18462 44952 18523 45006
rect 19198 44975 19258 45152
rect 19198 44952 19259 44975
rect 14043 44172 14103 44952
rect 16987 44588 17047 44952
rect 17721 44591 17781 44952
rect 16968 44579 17072 44588
rect 16968 44509 16982 44579
rect 17052 44509 17072 44579
rect 16968 44491 17072 44509
rect 17700 44580 17804 44591
rect 17700 44510 17716 44580
rect 17786 44510 17804 44580
rect 17700 44494 17804 44510
rect 14040 44171 14106 44172
rect 13312 44163 13378 44164
rect 13312 44099 13313 44163
rect 13377 44099 13378 44163
rect 14040 44107 14041 44171
rect 14105 44107 14106 44171
rect 14040 44106 14106 44107
rect 13312 44098 13378 44099
rect 12555 42728 12671 42734
rect 12555 42664 12581 42728
rect 12645 42664 12671 42728
rect 12555 42647 12671 42664
rect 18463 42186 18523 44952
rect 9800 29585 9878 29691
rect 9984 29585 10100 29691
rect 9263 24447 9424 24485
rect 9263 24377 9308 24447
rect 9378 24377 9424 24447
rect 9263 24325 9424 24377
rect 8862 17859 9023 17903
rect 8862 17789 8912 17859
rect 8982 17789 9023 17859
rect 8862 17743 9023 17789
rect 9800 17862 10100 29585
rect 9800 17722 9870 17862
rect 10002 17722 10100 17862
rect 9800 14044 10100 17722
rect 10565 42126 18523 42186
rect 9798 13936 10102 14044
rect 9798 13778 9894 13936
rect 10018 13778 10102 13936
rect 9798 13688 10102 13778
rect 5737 11909 5862 11921
rect 5737 11893 5756 11909
rect 842 11839 5756 11893
rect 5838 11839 5862 11909
rect 842 11831 5862 11839
rect 5737 11819 5862 11831
rect 6798 11915 6978 11945
rect 6798 11845 6844 11915
rect 6934 11845 6978 11915
rect 5738 11818 5861 11819
rect 4546 11454 4796 11488
rect 2672 11436 4796 11454
rect 2672 11320 4636 11436
rect 4726 11320 4796 11436
rect 2672 11274 4796 11320
rect 199 7231 501 7258
rect 199 7059 256 7231
rect 444 7059 501 7231
rect 199 7027 501 7059
rect 200 5098 500 7027
rect 200 4934 502 5098
rect 200 4762 256 4934
rect 444 4762 502 4934
rect 200 4634 502 4762
rect 200 1000 500 4634
rect 2672 1544 2852 11274
rect 4546 11272 4796 11274
rect 4612 10034 5152 10100
rect 4612 9786 4726 10034
rect 5044 9786 5152 10034
rect 4612 9712 5152 9786
rect 2674 1242 2852 1544
rect 4786 1496 4966 9712
rect 4785 1454 4966 1496
rect 4785 1383 4836 1454
rect 4910 1383 4966 1454
rect 4785 1348 4966 1383
rect 2674 1177 2737 1242
rect 2801 1177 2852 1242
rect 2674 1154 2852 1177
rect 6798 712 6978 11845
rect 9800 3546 10100 13688
rect 10565 12982 10625 42126
rect 19199 41942 19259 44952
rect 10830 41882 19259 41942
rect 10830 13130 10890 41882
rect 19934 41755 19994 45152
rect 10992 41695 19994 41755
rect 10992 13280 11052 41695
rect 20670 41596 20730 45152
rect 21406 44988 21466 45152
rect 11164 41536 20730 41596
rect 21402 44952 21466 44988
rect 22142 44970 22202 45152
rect 22878 44988 22938 45152
rect 22140 44952 22202 44970
rect 22877 44952 22938 44988
rect 23614 45042 23674 45152
rect 23614 44952 23675 45042
rect 24350 44992 24410 45152
rect 11164 13444 11224 41536
rect 21402 41396 21462 44952
rect 11328 41336 21462 41396
rect 11328 13590 11388 41336
rect 22140 41227 22200 44952
rect 11524 41167 22200 41227
rect 11524 13772 11584 41167
rect 22877 41041 22937 44952
rect 11742 40981 22937 41041
rect 11742 13913 11802 40981
rect 23615 40845 23675 44952
rect 11947 40785 23675 40845
rect 24348 44952 24410 44992
rect 11947 14068 12007 40785
rect 24348 40608 24408 44952
rect 12202 40548 24408 40608
rect 12202 14241 12262 40548
rect 25086 39552 25146 45152
rect 25822 45083 25882 45152
rect 13467 39492 25146 39552
rect 13467 37872 13527 39492
rect 25789 37927 25909 45083
rect 26558 45072 26618 45152
rect 27294 45080 27354 45152
rect 25788 37926 25910 37927
rect 13464 37871 13530 37872
rect 13464 37807 13465 37871
rect 13529 37807 13530 37871
rect 13464 37806 13530 37807
rect 25788 37806 25789 37926
rect 25909 37806 25910 37926
rect 25788 37805 25910 37806
rect 26508 30855 26628 45072
rect 27264 43154 27384 45080
rect 28030 45072 28090 45152
rect 27996 43488 28116 45072
rect 28766 45068 28826 45152
rect 28732 43924 28852 45068
rect 29502 45053 29562 45152
rect 30238 45117 30298 45152
rect 29470 44291 29590 45053
rect 30238 44952 30532 45117
rect 29464 44290 29596 44291
rect 29464 44170 29465 44290
rect 29595 44170 29596 44290
rect 29464 44169 29596 44170
rect 28721 43917 28865 43924
rect 28721 43787 28727 43917
rect 28857 43787 28865 43917
rect 28721 43781 28865 43787
rect 27984 43481 28128 43488
rect 27984 43351 27991 43481
rect 28121 43351 28128 43481
rect 27984 43345 28128 43351
rect 27253 43148 27397 43154
rect 27253 43018 27259 43148
rect 27389 43018 27397 43148
rect 27253 43011 27397 43018
rect 26507 30854 26629 30855
rect 26507 30734 26508 30854
rect 26628 30734 26629 30854
rect 26507 30733 26629 30734
rect 16187 28007 16367 28015
rect 16039 27993 16367 28007
rect 16039 27815 16056 27993
rect 16234 27815 16367 27993
rect 16039 27790 16367 27815
rect 15718 25063 16086 25137
rect 15718 24901 15803 25063
rect 15995 24901 16086 25063
rect 15718 24810 16086 24901
rect 12202 14181 14329 14241
rect 11947 14008 14037 14068
rect 11742 13853 13796 13913
rect 11524 13712 13605 13772
rect 11328 13530 13414 13590
rect 11164 13384 13209 13444
rect 10992 13220 13012 13280
rect 10830 13070 12812 13130
rect 10565 12922 12568 12982
rect 9800 3363 9875 3546
rect 10044 3363 10100 3546
rect 9800 1000 10100 3363
rect 10626 12321 10806 12355
rect 10626 12245 10679 12321
rect 10752 12245 10806 12321
rect 10626 1735 10806 12245
rect 11078 11469 11258 11501
rect 11078 11372 11131 11469
rect 11218 11372 11258 11469
rect 10625 1692 10807 1735
rect 10625 1601 10667 1692
rect 10761 1601 10807 1692
rect 10625 1556 10807 1601
rect 6798 532 9382 712
rect 370 0 550 200
rect 4786 0 4966 202
rect 9202 0 9382 532
rect 10626 374 10806 1556
rect 11078 775 11258 11372
rect 12508 1900 12568 12922
rect 12752 2054 12812 13070
rect 12952 2267 13012 13220
rect 13149 2420 13209 13384
rect 13354 2577 13414 13530
rect 13545 2696 13605 13712
rect 13736 2830 13796 13853
rect 13977 3009 14037 14008
rect 14269 3203 14329 14181
rect 14230 3138 14391 3203
rect 14230 3068 14264 3138
rect 14334 3068 14391 3138
rect 14230 3043 14391 3068
rect 13954 2997 14058 3009
rect 13954 2927 13972 2997
rect 14042 2927 14058 2997
rect 13954 2912 14058 2927
rect 13715 2815 13819 2830
rect 13715 2745 13731 2815
rect 13801 2745 13819 2815
rect 13715 2733 13819 2745
rect 13522 2683 13626 2696
rect 13522 2613 13540 2683
rect 13610 2613 13626 2683
rect 13522 2599 13626 2613
rect 13331 2565 13435 2577
rect 13331 2495 13349 2565
rect 13419 2495 13435 2565
rect 13331 2480 13435 2495
rect 13125 2405 13229 2420
rect 13125 2335 13144 2405
rect 13214 2335 13229 2405
rect 13125 2323 13229 2335
rect 12930 2256 13034 2267
rect 12930 2186 12947 2256
rect 13017 2186 13034 2256
rect 12930 2170 13034 2186
rect 12728 2041 12832 2054
rect 12728 1971 12747 2041
rect 12817 1971 12832 2041
rect 12728 1957 12832 1971
rect 12488 1887 12592 1900
rect 12488 1817 12503 1887
rect 12573 1817 12592 1887
rect 12488 1803 12592 1817
rect 15810 910 15990 24810
rect 16187 1296 16367 27790
rect 16592 27964 22216 27990
rect 16592 27852 22075 27964
rect 22177 27852 22216 27964
rect 16592 27810 22216 27852
rect 16592 1683 16772 27810
rect 30412 27176 30532 44952
rect 30974 44809 31034 45152
rect 31710 44952 31770 45152
rect 30856 44763 31216 44809
rect 30856 44626 30956 44763
rect 31070 44626 31216 44763
rect 30856 44549 31216 44626
rect 31445 44284 31565 44285
rect 31445 44166 31446 44284
rect 31564 44166 31565 44284
rect 31193 43911 31323 43918
rect 31193 43793 31197 43911
rect 31315 43793 31323 43911
rect 31193 43787 31323 43793
rect 30721 43476 30851 43481
rect 30721 43475 31102 43476
rect 30721 43357 30726 43475
rect 30844 43357 31102 43475
rect 30721 43356 31102 43357
rect 30721 43350 30851 43356
rect 30768 43142 30898 43149
rect 30768 43024 30774 43142
rect 30892 43024 30898 43142
rect 30768 43018 30898 43024
rect 30406 27175 30538 27176
rect 30406 27055 30407 27175
rect 30537 27055 30538 27175
rect 30406 27054 30538 27055
rect 30773 17917 30893 43018
rect 30772 17916 30894 17917
rect 30772 17796 30773 17916
rect 30893 17796 30894 17916
rect 30772 17795 30894 17796
rect 30982 13837 31102 43356
rect 30981 13836 31103 13837
rect 30981 13716 30982 13836
rect 31102 13716 31103 13836
rect 30981 13715 31103 13716
rect 31196 9757 31316 43787
rect 31195 9756 31317 9757
rect 31195 9636 31196 9756
rect 31316 9636 31317 9756
rect 31195 9635 31317 9636
rect 31445 5683 31565 44166
rect 31440 5676 31571 5683
rect 31440 5556 31445 5676
rect 31565 5556 31571 5676
rect 31440 5550 31571 5556
rect 16592 1636 31462 1683
rect 16592 1552 16642 1636
rect 16729 1552 31462 1636
rect 16592 1503 31462 1552
rect 16187 1243 27046 1296
rect 16187 1151 16248 1243
rect 16346 1151 27046 1243
rect 16187 1116 27046 1151
rect 11078 595 15194 775
rect 15810 730 22630 910
rect 15014 486 15194 595
rect 10626 194 13798 374
rect 15014 306 18214 486
rect 13618 0 13798 194
rect 18034 0 18214 306
rect 22450 0 22630 730
rect 26866 0 27046 1116
rect 31282 0 31462 1503
use mux_inv_demux_buff_comp  mux_inv_demux_buff_comp_0
timestamp 1717183646
transform 1 0 7640 0 1 26527
box -6162 -20493 1060 5158
use pwm_generator  pwm_generator_0
timestamp 1717180972
transform 1 0 17108 0 1 3644
box 0 0 14457 16601
use sky130_fd_pr__res_xhigh_po_0p35_NM7GYR  sky130_fd_pr__res_xhigh_po_0p35_NM7GYR_0
timestamp 1717180972
transform 1 0 1239 0 1 3856
box -35 -532 35 532
use Top  Top_0
timestamp 1717180972
transform 1 0 13146 0 1 27462
box 0 0 11954 14098
use vo2  vo2_0
timestamp 1717180972
transform 1 0 11460 0 1 4322
box 350 -2768 424 2611
use voltagedivider  voltagedivider_0
timestamp 1717180972
transform 1 0 1000 0 1 7708
box 205 -1952 276 4058
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
