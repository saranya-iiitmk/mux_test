magic
tech sky130B
magscale 1 2
timestamp 1717174014
<< xpolycontact >>
rect -35 600 35 1032
rect -35 -1032 35 -600
<< xpolyres >>
rect -35 -600 35 600
<< viali >>
rect -19 617 19 1014
rect -19 -1014 19 -617
<< metal1 >>
rect -25 1014 25 1026
rect -25 617 -19 1014
rect 19 617 25 1014
rect -25 605 25 617
rect -25 -617 25 -605
rect -25 -1014 -19 -617
rect 19 -1014 25 -617
rect -25 -1026 25 -1014
<< res0p35 >>
rect -37 -602 37 602
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 6.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 35.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
