magic
tech sky130A
timestamp 1717137789
<< error_s >>
rect 0 226 153 388
rect 18 62 47 162
rect 62 62 91 162
rect 106 62 135 162
<< poly >>
rect 47 212 62 247
rect 47 197 106 212
rect 91 175 106 197
use mux_unitcell  mux_unitcell_0
timestamp 1717137789
transform 1 0 364 0 1 -45
box -364 94 -255 433
use mux_unitcell  mux_unitcell_1
timestamp 1717137789
transform -1 0 -211 0 1 -45
box -364 94 -255 433
<< end >>
