magic
tech sky130A
magscale 1 2
timestamp 1717183646
<< nwell >>
rect -1290 -13139 -1256 -13076
rect -910 -13207 -741 -12810
rect -1290 -13357 -1256 -13323
<< psubdiff >>
rect -824 -12613 -678 -12560
rect -824 -12707 -787 -12613
rect -718 -12707 -678 -12613
rect -824 -12750 -678 -12707
<< nsubdiff >>
rect -889 -12980 -789 -12954
rect -889 -13030 -866 -12980
rect -813 -13030 -789 -12980
rect -889 -13057 -789 -13030
<< psubdiffcont >>
rect -787 -12707 -718 -12613
<< nsubdiffcont >>
rect -866 -13030 -813 -12980
<< poly >>
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -2160 -12611 -2023 -12586
rect -2109 -12768 -2078 -12611
rect -2328 -12800 -2078 -12768
rect -2260 -13575 -2051 -13545
rect -2081 -13771 -2051 -13575
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -2130 -13882 -1992 -13859
<< polycont >>
rect -2126 -12586 -2059 -12521
rect -2094 -13859 -2027 -13794
<< locali >>
rect -4672 3115 -4337 3183
rect -4672 2991 -4591 3115
rect -4444 3073 -4337 3115
rect -4444 3039 -3946 3073
rect -4444 2991 -4337 3039
rect -4672 2928 -4337 2991
rect -4794 -4600 -4491 -4530
rect -4794 -4714 -4710 -4600
rect -4584 -4636 -4491 -4600
rect -4584 -4670 -3990 -4636
rect -4584 -4714 -4491 -4670
rect -4794 -4783 -4491 -4714
rect -788 -12448 -714 -12437
rect -788 -12483 -764 -12448
rect -730 -12483 -714 -12448
rect -788 -12499 -714 -12483
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -778 -12560 -723 -12499
rect -2160 -12611 -2023 -12586
rect -824 -12613 -678 -12560
rect -1433 -12644 -1359 -12628
rect -1433 -12679 -1412 -12644
rect -1378 -12679 -1359 -12644
rect -824 -12647 -787 -12613
rect -1433 -12696 -1359 -12679
rect -923 -12681 -787 -12647
rect -824 -12707 -787 -12681
rect -718 -12636 -678 -12613
rect -718 -12670 -551 -12636
rect -718 -12707 -678 -12670
rect -824 -12750 -678 -12707
rect -889 -12980 -789 -12954
rect -889 -12985 -866 -12980
rect -928 -13021 -866 -12985
rect -889 -13030 -866 -13021
rect -813 -13030 -789 -12980
rect -889 -13057 -789 -13030
rect -3642 -13081 -3540 -13065
rect -3642 -13121 -3615 -13081
rect -3574 -13082 -3540 -13081
rect -3574 -13121 -3423 -13082
rect -3642 -13124 -3423 -13121
rect -3642 -13139 -3540 -13124
rect -1290 -13140 -1256 -13076
rect -852 -13130 -818 -13057
rect -1307 -13152 -1239 -13140
rect -1307 -13186 -1291 -13152
rect -1257 -13186 -1239 -13152
rect -1307 -13195 -1239 -13186
rect -872 -13145 -790 -13130
rect -872 -13185 -847 -13145
rect -810 -13185 -790 -13145
rect -1290 -13357 -1256 -13195
rect -872 -13196 -790 -13185
rect -852 -13357 -818 -13196
rect -585 -13332 -551 -12670
rect -613 -13342 -522 -13332
rect -613 -13394 -595 -13342
rect -541 -13394 -522 -13342
rect -613 -13408 -522 -13394
rect -3757 -13632 -3234 -13630
rect -3826 -13673 -3234 -13632
rect -585 -13661 -551 -13408
rect -3826 -13675 -3303 -13673
rect -3826 -13783 -3757 -13675
rect -3854 -13870 -3730 -13783
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -2130 -13882 -1992 -13859
rect -1299 -14066 -1265 -13661
rect -845 -13695 -551 -13661
rect -585 -14066 -551 -13695
rect -1299 -14100 -551 -14066
<< viali >>
rect -4591 2991 -4444 3115
rect -4710 -4714 -4584 -4600
rect -764 -12483 -730 -12448
rect -2126 -12586 -2059 -12521
rect -1412 -12679 -1378 -12644
rect -3615 -13121 -3574 -13081
rect -1291 -13186 -1257 -13152
rect -847 -13185 -810 -13145
rect -595 -13394 -541 -13342
rect -2094 -13859 -2027 -13794
<< metal1 >>
rect -4672 3115 -4337 3183
rect -4672 2991 -4591 3115
rect -4444 2991 -4337 3115
rect -4672 2928 -4337 2991
rect -5507 1688 -4164 1722
rect -5507 -5674 -5473 1688
rect -4198 1108 -4164 1688
rect -4794 -4600 -4491 -4530
rect -4794 -4714 -4710 -4600
rect -4584 -4714 -4491 -4600
rect -4794 -4783 -4491 -4714
rect -5507 -5708 -4208 -5674
rect -4242 -6497 -4208 -5708
rect -6162 -11922 -5989 -11903
rect -6162 -11983 -6125 -11922
rect -6043 -11937 -5989 -11922
rect -6043 -11971 -496 -11937
rect -6043 -11983 -5989 -11971
rect -6162 -12011 -5989 -11983
rect -788 -12448 -714 -12437
rect -788 -12453 -764 -12448
rect -1407 -12482 -764 -12453
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -2160 -12611 -2023 -12586
rect -1407 -12628 -1378 -12482
rect -788 -12483 -764 -12482
rect -730 -12483 -714 -12448
rect -788 -12499 -714 -12483
rect -1433 -12644 -1359 -12628
rect -1433 -12679 -1412 -12644
rect -1378 -12679 -1359 -12644
rect -1433 -12696 -1359 -12679
rect -6160 -12732 -5990 -12696
rect -6160 -12808 -6112 -12732
rect -6053 -12759 -5990 -12732
rect -6053 -12808 -3564 -12759
rect -6160 -12848 -5990 -12808
rect -3613 -13065 -3564 -12808
rect -3642 -13081 -3540 -13065
rect -3642 -13121 -3615 -13081
rect -3574 -13121 -3540 -13081
rect -3642 -13139 -3540 -13121
rect -1307 -13150 -1239 -13140
rect -872 -13145 -790 -13130
rect -872 -13150 -847 -13145
rect -1307 -13152 -847 -13150
rect -1307 -13186 -1291 -13152
rect -1257 -13185 -847 -13152
rect -810 -13146 -790 -13145
rect -530 -13146 -496 -11971
rect -810 -13180 -496 -13146
rect -810 -13185 -790 -13180
rect -1257 -13186 -1239 -13185
rect -1307 -13195 -1239 -13186
rect -872 -13196 -790 -13185
rect -613 -13342 -522 -13332
rect -613 -13394 -595 -13342
rect -541 -13394 -522 -13342
rect -613 -13408 -522 -13394
rect -3854 -13870 -3730 -13783
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -2130 -13882 -1992 -13859
<< via1 >>
rect -4591 2991 -4444 3115
rect -4710 -4714 -4584 -4600
rect -6125 -11983 -6043 -11922
rect -2126 -12586 -2059 -12521
rect -6112 -12808 -6053 -12732
rect -595 -13394 -541 -13342
rect -2094 -13859 -2027 -13794
<< metal2 >>
rect -6161 3084 -5989 5158
rect -4672 3115 -4337 3183
rect -4672 3084 -4591 3115
rect -6161 3002 -4591 3084
rect -6161 -4605 -5989 3002
rect -4672 2991 -4591 3002
rect -4444 2991 -4337 3115
rect -4672 2928 -4337 2991
rect -4794 -4600 -4491 -4530
rect -4794 -4605 -4710 -4600
rect -6161 -4710 -4710 -4605
rect -6161 -11903 -5989 -4710
rect -4794 -4714 -4710 -4710
rect -4584 -4714 -4491 -4600
rect -4794 -4783 -4491 -4714
rect 885 -11251 1058 -10659
rect 883 -11302 1058 -11251
rect 883 -11372 931 -11302
rect 1010 -11372 1058 -11302
rect 883 -11418 1058 -11372
rect -6162 -11922 -5989 -11903
rect -6162 -11983 -6125 -11922
rect -6043 -11983 -5989 -11922
rect -6162 -12011 -5989 -11983
rect -6161 -12732 -5989 -12011
rect 885 -11697 1058 -11418
rect 885 -11761 1060 -11697
rect 885 -11831 932 -11761
rect 1011 -11831 1060 -11761
rect 885 -11904 1060 -11831
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -2160 -12611 -2023 -12586
rect -6161 -12808 -6112 -12732
rect -6053 -12808 -5989 -12732
rect -6161 -15321 -5989 -12808
rect -613 -13341 -522 -13332
rect 885 -13341 1058 -11904
rect -613 -13342 1058 -13341
rect -613 -13394 -595 -13342
rect -541 -13393 1058 -13342
rect -541 -13394 -522 -13393
rect -613 -13408 -522 -13394
rect -3854 -13870 -3730 -13783
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -3826 -14440 -3757 -13870
rect -2130 -13882 -1992 -13859
rect 885 -14440 1058 -13393
rect -3826 -14509 1058 -14440
rect 885 -15321 1058 -14509
rect 885 -20493 1058 -20369
<< via2 >>
rect 931 -11372 1010 -11302
rect 932 -11831 1011 -11761
rect -2126 -12586 -2059 -12521
rect -2094 -13859 -2027 -13794
<< metal3 >>
rect -786 -1956 -702 -1581
rect -786 -2040 499 -1956
rect -844 -11771 -768 -9183
rect 385 -11285 469 -2040
rect 883 -11285 1058 -11251
rect 385 -11302 1058 -11285
rect 385 -11369 931 -11302
rect 883 -11372 931 -11369
rect 1010 -11372 1058 -11302
rect 883 -11418 1058 -11372
rect 885 -11761 1060 -11697
rect 885 -11771 932 -11761
rect -844 -11831 932 -11771
rect 1011 -11831 1060 -11761
rect -844 -11847 1060 -11831
rect 885 -11904 1060 -11847
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -2160 -12611 -2023 -12586
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -2130 -13882 -1992 -13859
<< via3 >>
rect -2126 -12586 -2059 -12521
rect -2094 -13859 -2027 -13794
<< metal4 >>
rect -5815 4939 -985 5043
rect -5815 -11683 -5711 4939
rect -1089 4760 -985 4939
rect -1090 4698 -985 4760
rect -1089 4656 -985 4698
rect -1133 -2443 182 -2339
rect -1133 -2952 -1029 -2443
rect -5815 -11787 -2048 -11683
rect -2133 -12499 -2048 -11787
rect -2160 -12521 -2023 -12499
rect -2160 -12586 -2126 -12521
rect -2059 -12586 -2023 -12521
rect -2160 -12611 -2023 -12586
rect -2130 -13794 -1992 -13771
rect -2130 -13859 -2094 -13794
rect -2027 -13859 -1992 -13794
rect -2130 -13882 -1992 -13859
rect -2110 -14086 -2005 -13882
rect -2110 -14238 -2004 -14086
rect 78 -14238 182 -2443
rect -2110 -14342 182 -14238
use comparator  comparator_0
timestamp 1717183646
transform 1 0 -10006 0 1 6500
box 4736 -8254 9501 -1774
use comparator  comparator_1
timestamp 1717183646
transform 1 0 -10050 0 1 -1094
box 4736 -8254 9501 -1774
use mux_inv_demux_buff  mux_inv_demux_buff_1
timestamp 1717180972
transform 1 0 -2980 0 1 -13873
box -890 -424 2169 1662
<< labels >>
rlabel metal2 912 -15293 1035 -15093 1 GND
rlabel metal2 -6137 -15180 -6014 -14980 1 VDD
<< end >>
