VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mixed_signal_pulse_gen
  CLASS BLOCK ;
  FOREIGN tt_um_mixed_signal_pulse_gen ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.704000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.796500 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.096500 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.722900 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 1.085200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 71.060 193.015 119.740 194.620 ;
      LAYER pwell ;
        RECT 71.255 191.815 72.625 192.625 ;
        RECT 72.635 191.815 78.145 192.625 ;
        RECT 78.155 191.815 80.905 192.625 ;
        RECT 80.915 191.815 83.655 192.495 ;
        RECT 84.145 191.900 84.575 192.685 ;
        RECT 84.595 191.815 85.965 192.625 ;
        RECT 86.070 192.495 86.990 192.725 ;
        RECT 86.070 191.815 89.535 192.495 ;
        RECT 89.655 191.815 95.165 192.625 ;
        RECT 95.175 191.815 97.005 192.625 ;
        RECT 97.025 191.900 97.455 192.685 ;
        RECT 97.475 191.815 100.225 192.625 ;
        RECT 101.285 192.495 102.215 192.725 ;
        RECT 100.380 191.815 102.215 192.495 ;
        RECT 102.535 191.815 108.045 192.625 ;
        RECT 108.055 191.815 109.885 192.625 ;
        RECT 109.905 191.900 110.335 192.685 ;
        RECT 110.815 191.815 113.555 192.495 ;
        RECT 113.575 191.815 117.245 192.625 ;
        RECT 118.175 191.815 119.545 192.625 ;
        RECT 71.395 191.605 71.565 191.815 ;
        RECT 72.775 191.605 72.945 191.815 ;
        RECT 74.155 191.605 74.325 191.795 ;
        RECT 76.910 191.655 77.030 191.765 ;
        RECT 78.295 191.625 78.465 191.815 ;
        RECT 81.055 191.625 81.225 191.815 ;
        RECT 82.430 191.605 82.600 191.795 ;
        RECT 82.890 191.605 83.060 191.795 ;
        RECT 83.810 191.655 83.930 191.765 ;
        RECT 84.275 191.605 84.445 191.795 ;
        RECT 84.735 191.625 84.905 191.815 ;
        RECT 89.335 191.625 89.505 191.815 ;
        RECT 89.795 191.625 89.965 191.815 ;
        RECT 93.935 191.605 94.105 191.795 ;
        RECT 95.315 191.625 95.485 191.815 ;
        RECT 95.770 191.605 95.940 191.795 ;
        RECT 96.245 191.650 96.405 191.760 ;
        RECT 97.615 191.625 97.785 191.815 ;
        RECT 100.380 191.795 100.545 191.815 ;
        RECT 100.375 191.625 100.545 191.795 ;
        RECT 100.835 191.605 101.005 191.795 ;
        RECT 101.295 191.605 101.465 191.795 ;
        RECT 102.675 191.625 102.845 191.815 ;
        RECT 104.055 191.605 104.225 191.795 ;
        RECT 105.900 191.605 106.070 191.795 ;
        RECT 108.195 191.625 108.365 191.815 ;
        RECT 110.490 191.655 110.610 191.765 ;
        RECT 110.955 191.625 111.125 191.815 ;
        RECT 111.415 191.605 111.585 191.795 ;
        RECT 113.715 191.625 113.885 191.815 ;
        RECT 117.405 191.660 117.565 191.770 ;
        RECT 117.845 191.605 118.015 191.795 ;
        RECT 119.235 191.605 119.405 191.815 ;
        RECT 71.255 190.795 72.625 191.605 ;
        RECT 72.635 190.825 74.005 191.605 ;
        RECT 74.015 190.795 76.765 191.605 ;
        RECT 77.235 190.925 82.745 191.605 ;
        RECT 77.235 190.695 78.625 190.925 ;
        RECT 82.775 190.695 84.125 191.605 ;
        RECT 84.135 190.795 86.885 191.605 ;
        RECT 86.935 190.925 94.245 191.605 ;
        RECT 86.935 190.695 88.285 190.925 ;
        RECT 89.820 190.705 90.730 190.925 ;
        RECT 94.255 190.695 96.085 191.605 ;
        RECT 97.025 190.735 97.455 191.520 ;
        RECT 97.570 190.925 101.035 191.605 ;
        RECT 97.570 190.695 98.490 190.925 ;
        RECT 101.165 190.695 103.895 191.605 ;
        RECT 103.915 190.795 105.745 191.605 ;
        RECT 105.755 190.925 111.265 191.605 ;
        RECT 109.875 190.695 111.265 190.925 ;
        RECT 111.275 190.795 116.785 191.605 ;
        RECT 116.795 190.825 118.165 191.605 ;
        RECT 118.175 190.795 119.545 191.605 ;
      LAYER nwell ;
        RECT 71.060 187.575 119.740 190.405 ;
      LAYER pwell ;
        RECT 71.255 186.375 72.625 187.185 ;
        RECT 72.635 186.375 78.145 187.185 ;
        RECT 78.155 186.375 79.985 187.185 ;
        RECT 83.175 187.085 84.125 187.285 ;
        RECT 80.455 186.405 84.125 187.085 ;
        RECT 84.145 186.460 84.575 187.245 ;
        RECT 88.110 187.055 89.020 187.275 ;
        RECT 90.555 187.055 91.905 187.285 ;
        RECT 71.395 186.165 71.565 186.375 ;
        RECT 72.775 186.165 72.945 186.375 ;
        RECT 78.295 186.165 78.465 186.375 ;
        RECT 80.130 186.215 80.250 186.325 ;
        RECT 80.600 186.185 80.770 186.405 ;
        RECT 83.175 186.375 84.125 186.405 ;
        RECT 84.595 186.375 91.905 187.055 ;
        RECT 92.050 187.055 92.970 187.285 ;
        RECT 92.050 186.375 95.515 187.055 ;
        RECT 95.645 186.375 96.995 187.285 ;
        RECT 100.530 187.055 101.440 187.275 ;
        RECT 102.975 187.055 104.325 187.285 ;
        RECT 97.015 186.375 104.325 187.055 ;
        RECT 104.455 186.375 107.455 187.285 ;
        RECT 107.595 186.375 108.945 187.285 ;
        RECT 109.905 186.460 110.335 187.245 ;
        RECT 113.080 187.085 114.025 187.285 ;
        RECT 111.275 186.405 114.025 187.085 ;
        RECT 84.735 186.185 84.905 186.375 ;
        RECT 71.255 185.355 72.625 186.165 ;
        RECT 72.635 185.355 78.145 186.165 ;
        RECT 78.155 185.355 83.665 186.165 ;
        RECT 83.675 186.135 84.620 186.165 ;
        RECT 86.575 186.135 86.745 186.355 ;
        RECT 91.200 186.185 91.370 186.355 ;
        RECT 91.200 186.165 91.310 186.185 ;
        RECT 91.635 186.165 91.805 186.355 ;
        RECT 93.475 186.165 93.645 186.355 ;
        RECT 95.315 186.185 95.485 186.375 ;
        RECT 95.775 186.185 95.945 186.375 ;
        RECT 97.155 186.185 97.325 186.375 ;
        RECT 97.625 186.210 97.785 186.320 ;
        RECT 98.540 186.165 98.710 186.355 ;
        RECT 83.675 185.935 86.745 186.135 ;
        RECT 83.675 185.455 86.885 185.935 ;
        RECT 83.675 185.255 84.620 185.455 ;
        RECT 85.955 185.255 86.885 185.455 ;
        RECT 86.895 185.485 91.310 186.165 ;
        RECT 86.895 185.255 90.825 185.485 ;
        RECT 91.495 185.355 93.325 186.165 ;
        RECT 93.445 185.485 96.910 186.165 ;
        RECT 95.990 185.255 96.910 185.485 ;
        RECT 97.025 185.295 97.455 186.080 ;
        RECT 98.395 185.485 102.065 186.165 ;
        RECT 102.210 186.135 102.380 186.355 ;
        RECT 104.515 186.165 104.685 186.375 ;
        RECT 107.275 186.165 107.445 186.355 ;
        RECT 107.740 186.185 107.910 186.375 ;
        RECT 108.655 186.165 108.825 186.355 ;
        RECT 109.115 186.165 109.285 186.355 ;
        RECT 110.505 186.220 110.665 186.330 ;
        RECT 110.955 186.165 111.125 186.355 ;
        RECT 111.420 186.185 111.590 186.405 ;
        RECT 113.080 186.375 114.025 186.405 ;
        RECT 114.035 186.375 115.405 187.155 ;
        RECT 115.415 186.375 118.165 187.185 ;
        RECT 118.175 186.375 119.545 187.185 ;
        RECT 115.095 186.185 115.265 186.375 ;
        RECT 115.555 186.185 115.725 186.375 ;
        RECT 119.235 186.165 119.405 186.375 ;
        RECT 103.410 186.135 104.365 186.165 ;
        RECT 98.395 185.255 99.320 185.485 ;
        RECT 102.085 185.455 104.365 186.135 ;
        RECT 103.410 185.255 104.365 185.455 ;
        RECT 104.375 185.355 106.205 186.165 ;
        RECT 106.215 185.385 107.585 186.165 ;
        RECT 107.595 185.385 108.965 186.165 ;
        RECT 108.975 185.355 110.805 186.165 ;
        RECT 110.815 185.485 118.125 186.165 ;
        RECT 114.330 185.265 115.240 185.485 ;
        RECT 116.775 185.255 118.125 185.485 ;
        RECT 118.175 185.355 119.545 186.165 ;
      LAYER nwell ;
        RECT 71.060 182.135 119.740 184.965 ;
      LAYER pwell ;
        RECT 71.255 180.935 72.625 181.745 ;
        RECT 72.635 180.935 78.145 181.745 ;
        RECT 78.155 180.935 83.665 181.745 ;
        RECT 84.145 181.020 84.575 181.805 ;
        RECT 84.595 180.935 86.425 181.745 ;
        RECT 89.550 181.615 90.470 181.845 ;
        RECT 87.005 180.935 90.470 181.615 ;
        RECT 90.575 180.935 92.405 181.745 ;
        RECT 94.220 181.645 95.165 181.845 ;
        RECT 92.415 180.965 95.165 181.645 ;
        RECT 71.395 180.725 71.565 180.935 ;
        RECT 72.775 180.745 72.945 180.935 ;
        RECT 73.695 180.725 73.865 180.915 ;
        RECT 78.295 180.745 78.465 180.935 ;
        RECT 82.895 180.725 83.065 180.915 ;
        RECT 84.735 180.885 84.905 180.935 ;
        RECT 83.810 180.775 83.930 180.885 ;
        RECT 84.730 180.775 84.905 180.885 ;
        RECT 84.735 180.745 84.905 180.775 ;
        RECT 86.105 180.725 86.275 180.915 ;
        RECT 86.575 180.885 86.745 180.915 ;
        RECT 86.570 180.775 86.745 180.885 ;
        RECT 86.575 180.725 86.745 180.775 ;
        RECT 87.035 180.745 87.205 180.935 ;
        RECT 90.715 180.745 90.885 180.935 ;
        RECT 92.095 180.725 92.265 180.915 ;
        RECT 92.560 180.745 92.730 180.965 ;
        RECT 94.220 180.935 95.165 180.965 ;
        RECT 95.635 180.935 97.825 181.845 ;
        RECT 97.935 180.935 103.445 181.745 ;
        RECT 103.930 181.615 105.300 181.845 ;
        RECT 103.930 180.935 106.205 181.615 ;
        RECT 106.215 180.935 109.885 181.745 ;
        RECT 109.905 181.020 110.335 181.805 ;
        RECT 110.355 180.935 113.105 181.745 ;
        RECT 113.125 180.935 114.475 181.845 ;
        RECT 114.590 181.615 115.510 181.845 ;
        RECT 114.590 180.935 118.055 181.615 ;
        RECT 118.175 180.935 119.545 181.745 ;
        RECT 95.780 180.915 95.950 180.935 ;
        RECT 95.310 180.775 95.430 180.885 ;
        RECT 95.775 180.745 95.950 180.915 ;
        RECT 98.075 180.745 98.245 180.935 ;
        RECT 99.455 180.745 99.625 180.915 ;
        RECT 95.775 180.725 95.945 180.745 ;
        RECT 99.455 180.725 99.620 180.745 ;
        RECT 99.915 180.725 100.085 180.915 ;
        RECT 101.295 180.725 101.465 180.915 ;
        RECT 103.590 180.775 103.710 180.885 ;
        RECT 104.055 180.725 104.225 180.915 ;
        RECT 105.435 180.725 105.605 180.915 ;
        RECT 105.890 180.745 106.060 180.935 ;
        RECT 106.355 180.745 106.525 180.935 ;
        RECT 110.495 180.745 110.665 180.935 ;
        RECT 112.795 180.725 112.965 180.915 ;
        RECT 114.175 180.745 114.345 180.935 ;
        RECT 117.855 180.745 118.025 180.935 ;
        RECT 119.235 180.725 119.405 180.935 ;
        RECT 71.255 179.915 72.625 180.725 ;
        RECT 73.555 180.045 82.745 180.725 ;
        RECT 78.065 179.825 78.995 180.045 ;
        RECT 81.825 179.815 82.745 180.045 ;
        RECT 82.755 179.915 84.585 180.725 ;
        RECT 85.055 179.945 86.425 180.725 ;
        RECT 86.435 179.915 91.945 180.725 ;
        RECT 91.955 179.915 95.625 180.725 ;
        RECT 95.635 179.915 97.005 180.725 ;
        RECT 97.025 179.855 97.455 180.640 ;
        RECT 97.785 180.045 99.620 180.725 ;
        RECT 97.785 179.815 98.715 180.045 ;
        RECT 99.775 179.915 101.145 180.725 ;
        RECT 101.165 179.815 103.895 180.725 ;
        RECT 103.915 179.915 105.285 180.725 ;
        RECT 105.295 180.045 112.605 180.725 ;
        RECT 108.810 179.825 109.720 180.045 ;
        RECT 111.255 179.815 112.605 180.045 ;
        RECT 112.655 179.915 118.165 180.725 ;
        RECT 118.175 179.915 119.545 180.725 ;
      LAYER nwell ;
        RECT 71.060 176.695 119.740 179.525 ;
      LAYER pwell ;
        RECT 71.255 175.495 72.625 176.305 ;
        RECT 73.555 175.495 76.725 176.405 ;
        RECT 76.775 175.495 80.445 176.305 ;
        RECT 80.915 175.495 84.085 176.405 ;
        RECT 84.145 175.580 84.575 176.365 ;
        RECT 84.595 175.495 90.105 176.305 ;
        RECT 90.115 175.495 91.945 176.305 ;
        RECT 101.250 176.175 102.170 176.405 ;
        RECT 105.390 176.175 106.310 176.405 ;
        RECT 91.955 175.495 101.060 176.175 ;
        RECT 101.250 175.495 104.715 176.175 ;
        RECT 105.390 175.495 108.855 176.175 ;
        RECT 109.905 175.580 110.335 176.365 ;
        RECT 110.355 176.175 111.285 176.405 ;
        RECT 110.355 175.495 114.255 176.175 ;
        RECT 114.495 175.495 115.845 176.405 ;
        RECT 115.875 175.495 117.225 176.405 ;
        RECT 118.175 175.495 119.545 176.305 ;
        RECT 71.395 175.285 71.565 175.495 ;
        RECT 72.775 175.285 72.945 175.475 ;
        RECT 74.155 175.285 74.325 175.475 ;
        RECT 76.455 175.305 76.625 175.495 ;
        RECT 76.915 175.305 77.085 175.495 ;
        RECT 80.590 175.335 80.710 175.445 ;
        RECT 83.355 175.285 83.525 175.475 ;
        RECT 83.815 175.305 83.985 175.495 ;
        RECT 84.735 175.285 84.905 175.495 ;
        RECT 90.255 175.305 90.425 175.495 ;
        RECT 92.095 175.305 92.265 175.495 ;
        RECT 93.930 175.335 94.050 175.445 ;
        RECT 94.395 175.285 94.565 175.475 ;
        RECT 97.615 175.285 97.785 175.475 ;
        RECT 104.515 175.305 104.685 175.495 ;
        RECT 104.970 175.335 105.090 175.445 ;
        RECT 108.655 175.305 108.825 175.495 ;
        RECT 108.840 175.285 109.010 175.475 ;
        RECT 109.125 175.340 109.285 175.450 ;
        RECT 110.490 175.285 110.660 175.475 ;
        RECT 110.770 175.305 110.940 175.495 ;
        RECT 110.950 175.335 111.070 175.445 ;
        RECT 114.820 175.285 114.990 175.475 ;
        RECT 115.560 175.305 115.730 175.495 ;
        RECT 116.940 175.305 117.110 175.495 ;
        RECT 117.395 175.305 117.565 175.475 ;
        RECT 117.850 175.335 117.970 175.445 ;
        RECT 117.395 175.285 117.560 175.305 ;
        RECT 119.235 175.285 119.405 175.495 ;
        RECT 71.255 174.475 72.625 175.285 ;
        RECT 72.635 174.475 74.005 175.285 ;
        RECT 74.015 174.605 83.205 175.285 ;
        RECT 78.525 174.385 79.455 174.605 ;
        RECT 82.285 174.375 83.205 174.605 ;
        RECT 83.215 174.475 84.585 175.285 ;
        RECT 84.595 174.605 93.785 175.285 ;
        RECT 89.105 174.385 90.035 174.605 ;
        RECT 92.865 174.375 93.785 174.605 ;
        RECT 94.255 174.375 97.005 175.285 ;
        RECT 97.025 174.415 97.455 175.200 ;
        RECT 97.475 174.605 104.785 175.285 ;
        RECT 105.525 174.605 109.425 175.285 ;
        RECT 100.990 174.385 101.900 174.605 ;
        RECT 103.435 174.375 104.785 174.605 ;
        RECT 108.495 174.375 109.425 174.605 ;
        RECT 109.455 174.375 110.805 175.285 ;
        RECT 111.505 174.605 115.405 175.285 ;
        RECT 114.475 174.375 115.405 174.605 ;
        RECT 115.725 174.605 117.560 175.285 ;
        RECT 115.725 174.375 116.655 174.605 ;
        RECT 118.175 174.475 119.545 175.285 ;
      LAYER nwell ;
        RECT 71.060 171.255 119.740 174.085 ;
      LAYER pwell ;
        RECT 71.255 170.055 72.625 170.865 ;
        RECT 72.635 170.055 74.465 170.865 ;
        RECT 74.935 170.055 78.045 170.965 ;
        RECT 78.155 170.055 83.665 170.865 ;
        RECT 84.145 170.140 84.575 170.925 ;
        RECT 84.595 170.055 85.965 170.835 ;
        RECT 85.975 170.055 87.805 170.865 ;
        RECT 87.815 170.735 91.745 170.965 ;
        RECT 106.050 170.735 106.960 170.955 ;
        RECT 108.495 170.735 109.845 170.965 ;
        RECT 87.815 170.055 92.230 170.735 ;
        RECT 92.415 170.055 101.520 170.735 ;
        RECT 102.535 170.055 109.845 170.735 ;
        RECT 109.905 170.140 110.335 170.925 ;
        RECT 110.450 170.735 111.370 170.965 ;
        RECT 114.130 170.735 115.050 170.965 ;
        RECT 110.450 170.055 113.915 170.735 ;
        RECT 114.130 170.055 117.595 170.735 ;
        RECT 118.175 170.055 119.545 170.865 ;
        RECT 71.395 169.845 71.565 170.055 ;
        RECT 72.775 169.845 72.945 170.055 ;
        RECT 74.610 169.895 74.730 170.005 ;
        RECT 77.835 169.865 78.005 170.055 ;
        RECT 78.295 169.845 78.465 170.055 ;
        RECT 84.745 170.035 84.915 170.055 ;
        RECT 83.810 170.000 83.930 170.005 ;
        RECT 83.810 169.895 83.985 170.000 ;
        RECT 83.825 169.890 83.985 169.895 ;
        RECT 84.735 169.865 84.915 170.035 ;
        RECT 86.115 169.865 86.285 170.055 ;
        RECT 92.120 170.035 92.230 170.055 ;
        RECT 84.735 169.845 84.905 169.865 ;
        RECT 87.955 169.845 88.125 170.035 ;
        RECT 91.175 169.845 91.345 170.035 ;
        RECT 92.120 169.865 92.290 170.035 ;
        RECT 92.555 169.865 92.725 170.055 ;
        RECT 94.855 169.845 95.025 170.035 ;
        RECT 96.690 169.895 96.810 170.005 ;
        RECT 97.615 169.845 97.785 170.035 ;
        RECT 99.455 169.845 99.625 170.035 ;
        RECT 101.765 169.900 101.925 170.010 ;
        RECT 102.675 169.865 102.845 170.055 ;
        RECT 103.135 169.845 103.305 170.035 ;
        RECT 105.435 169.845 105.605 170.035 ;
        RECT 105.895 169.845 106.065 170.035 ;
        RECT 107.735 169.845 107.905 170.035 ;
        RECT 110.955 169.845 111.125 170.035 ;
        RECT 113.715 169.865 113.885 170.055 ;
        RECT 117.395 169.865 117.565 170.055 ;
        RECT 117.850 169.895 117.970 170.005 ;
        RECT 119.235 169.845 119.405 170.055 ;
        RECT 71.255 169.035 72.625 169.845 ;
        RECT 72.635 169.035 78.145 169.845 ;
        RECT 78.155 169.035 83.665 169.845 ;
        RECT 84.635 168.935 87.805 169.845 ;
        RECT 87.855 168.935 91.025 169.845 ;
        RECT 91.145 169.165 94.610 169.845 ;
        RECT 93.690 168.935 94.610 169.165 ;
        RECT 94.715 169.035 96.545 169.845 ;
        RECT 97.025 168.975 97.455 169.760 ;
        RECT 97.475 169.165 99.305 169.845 ;
        RECT 97.960 168.935 99.305 169.165 ;
        RECT 99.315 169.035 102.985 169.845 ;
        RECT 102.995 169.035 104.365 169.845 ;
        RECT 104.375 169.065 105.745 169.845 ;
        RECT 105.755 169.035 107.585 169.845 ;
        RECT 107.695 168.935 110.805 169.845 ;
        RECT 110.815 169.165 118.125 169.845 ;
        RECT 114.330 168.945 115.240 169.165 ;
        RECT 116.775 168.935 118.125 169.165 ;
        RECT 118.175 169.035 119.545 169.845 ;
      LAYER nwell ;
        RECT 71.060 165.815 119.740 168.645 ;
      LAYER pwell ;
        RECT 71.255 164.615 72.625 165.425 ;
        RECT 72.635 164.615 74.465 165.425 ;
        RECT 74.475 164.615 77.585 165.525 ;
        RECT 77.695 164.615 80.805 165.525 ;
        RECT 80.955 164.615 84.125 165.525 ;
        RECT 84.145 164.700 84.575 165.485 ;
        RECT 84.595 164.615 85.965 165.425 ;
        RECT 88.630 165.295 89.550 165.525 ;
        RECT 86.085 164.615 89.550 165.295 ;
        RECT 89.655 164.615 91.485 165.425 ;
        RECT 91.955 164.615 93.325 165.395 ;
        RECT 97.845 165.295 98.775 165.515 ;
        RECT 101.605 165.295 102.525 165.525 ;
        RECT 93.335 164.615 102.525 165.295 ;
        RECT 102.535 164.615 106.205 165.425 ;
        RECT 106.675 165.325 107.620 165.525 ;
        RECT 106.675 164.645 109.425 165.325 ;
        RECT 109.905 164.700 110.335 165.485 ;
        RECT 106.675 164.615 107.620 164.645 ;
        RECT 71.395 164.405 71.565 164.615 ;
        RECT 72.775 164.405 72.945 164.615 ;
        RECT 75.535 164.405 75.705 164.595 ;
        RECT 77.375 164.425 77.545 164.615 ;
        RECT 80.595 164.425 80.765 164.615 ;
        RECT 81.055 164.425 81.225 164.615 ;
        RECT 84.735 164.425 84.905 164.615 ;
        RECT 86.115 164.425 86.285 164.615 ;
        RECT 89.795 164.425 89.965 164.615 ;
        RECT 91.630 164.455 91.750 164.565 ;
        RECT 93.005 164.425 93.175 164.615 ;
        RECT 93.475 164.425 93.645 164.615 ;
        RECT 94.395 164.405 94.565 164.595 ;
        RECT 94.855 164.405 95.025 164.595 ;
        RECT 96.690 164.455 96.810 164.565 ;
        RECT 97.615 164.405 97.785 164.595 ;
        RECT 102.675 164.425 102.845 164.615 ;
        RECT 106.350 164.455 106.470 164.565 ;
        RECT 106.815 164.405 106.985 164.595 ;
        RECT 108.195 164.405 108.365 164.595 ;
        RECT 109.110 164.425 109.280 164.645 ;
        RECT 110.355 164.615 111.725 165.425 ;
        RECT 111.830 165.295 112.750 165.525 ;
        RECT 111.830 164.615 115.295 165.295 ;
        RECT 115.415 164.615 116.765 165.525 ;
        RECT 116.795 164.615 118.165 165.425 ;
        RECT 118.175 164.615 119.545 165.425 ;
        RECT 109.570 164.455 109.690 164.565 ;
        RECT 110.495 164.425 110.665 164.615 ;
        RECT 115.095 164.425 115.265 164.615 ;
        RECT 115.555 164.405 115.725 164.595 ;
        RECT 116.480 164.425 116.650 164.615 ;
        RECT 116.935 164.425 117.105 164.615 ;
        RECT 119.235 164.405 119.405 164.615 ;
        RECT 71.255 163.595 72.625 164.405 ;
        RECT 72.635 163.595 75.385 164.405 ;
        RECT 75.395 163.725 84.585 164.405 ;
        RECT 79.905 163.505 80.835 163.725 ;
        RECT 83.665 163.495 84.585 163.725 ;
        RECT 85.515 163.725 94.705 164.405 ;
        RECT 85.515 163.495 86.435 163.725 ;
        RECT 89.265 163.505 90.195 163.725 ;
        RECT 94.715 163.595 96.545 164.405 ;
        RECT 97.025 163.535 97.455 164.320 ;
        RECT 97.475 163.725 106.665 164.405 ;
        RECT 101.985 163.505 102.915 163.725 ;
        RECT 105.745 163.495 106.665 163.725 ;
        RECT 106.675 163.595 108.045 164.405 ;
        RECT 108.055 163.725 115.365 164.405 ;
        RECT 111.570 163.505 112.480 163.725 ;
        RECT 114.015 163.495 115.365 163.725 ;
        RECT 115.415 163.595 118.165 164.405 ;
        RECT 118.175 163.595 119.545 164.405 ;
      LAYER nwell ;
        RECT 71.060 160.375 119.740 163.205 ;
      LAYER pwell ;
        RECT 71.255 159.175 72.625 159.985 ;
        RECT 72.635 159.175 78.145 159.985 ;
        RECT 78.155 159.175 83.665 159.985 ;
        RECT 84.145 159.260 84.575 160.045 ;
        RECT 84.595 159.175 86.425 159.985 ;
        RECT 87.095 159.855 91.025 160.085 ;
        RECT 86.610 159.175 91.025 159.855 ;
        RECT 91.035 159.175 96.545 159.985 ;
        RECT 96.555 159.175 102.065 159.985 ;
        RECT 104.730 159.855 105.650 160.085 ;
        RECT 102.185 159.175 105.650 159.855 ;
        RECT 105.850 159.855 106.770 160.085 ;
        RECT 105.850 159.175 109.315 159.855 ;
        RECT 109.905 159.260 110.335 160.045 ;
        RECT 110.425 159.175 114.485 160.085 ;
        RECT 114.590 159.855 115.510 160.085 ;
        RECT 114.590 159.175 118.055 159.855 ;
        RECT 118.175 159.175 119.545 159.985 ;
        RECT 71.395 158.965 71.565 159.175 ;
        RECT 72.775 158.965 72.945 159.175 ;
        RECT 78.295 158.965 78.465 159.175 ;
        RECT 81.050 159.015 81.170 159.125 ;
        RECT 81.515 158.965 81.685 159.155 ;
        RECT 83.810 159.015 83.930 159.125 ;
        RECT 84.735 158.985 84.905 159.175 ;
        RECT 86.610 159.155 86.720 159.175 ;
        RECT 86.550 158.985 86.720 159.155 ;
        RECT 87.495 158.965 87.665 159.155 ;
        RECT 87.955 158.965 88.125 159.155 ;
        RECT 91.175 159.125 91.345 159.175 ;
        RECT 91.170 159.015 91.345 159.125 ;
        RECT 91.175 158.985 91.345 159.015 ;
        RECT 91.635 158.965 91.805 159.155 ;
        RECT 95.315 158.965 95.485 159.155 ;
        RECT 96.695 158.985 96.865 159.175 ;
        RECT 97.615 158.965 97.785 159.155 ;
        RECT 101.290 159.015 101.410 159.125 ;
        RECT 101.755 158.965 101.925 159.155 ;
        RECT 102.215 158.985 102.385 159.175 ;
        RECT 105.890 159.015 106.010 159.125 ;
        RECT 109.115 158.985 109.285 159.175 ;
        RECT 109.570 159.015 109.690 159.125 ;
        RECT 114.175 158.985 114.345 159.175 ;
        RECT 115.555 158.965 115.725 159.155 ;
        RECT 116.015 158.965 116.185 159.155 ;
        RECT 117.855 159.125 118.025 159.175 ;
        RECT 117.850 159.015 118.025 159.125 ;
        RECT 117.855 158.985 118.025 159.015 ;
        RECT 119.235 158.965 119.405 159.175 ;
        RECT 71.255 158.155 72.625 158.965 ;
        RECT 72.635 158.155 78.145 158.965 ;
        RECT 78.155 158.155 80.905 158.965 ;
        RECT 81.415 158.055 84.585 158.965 ;
        RECT 84.595 158.055 87.765 158.965 ;
        RECT 87.855 158.055 91.025 158.965 ;
        RECT 91.605 158.285 95.070 158.965 ;
        RECT 94.150 158.055 95.070 158.285 ;
        RECT 95.175 158.155 97.005 158.965 ;
        RECT 97.025 158.095 97.455 158.880 ;
        RECT 97.475 158.155 101.145 158.965 ;
        RECT 101.615 158.055 105.675 158.965 ;
        RECT 106.215 158.715 111.310 158.965 ;
        RECT 114.105 158.795 115.865 158.965 ;
        RECT 113.610 158.750 115.865 158.795 ;
        RECT 112.670 158.715 115.865 158.750 ;
        RECT 106.215 158.285 115.865 158.715 ;
        RECT 106.215 158.055 108.235 158.285 ;
        RECT 107.315 158.035 108.235 158.055 ;
        RECT 111.310 158.115 114.540 158.285 ;
        RECT 115.875 158.155 117.705 158.965 ;
        RECT 118.175 158.155 119.545 158.965 ;
        RECT 111.310 158.070 113.600 158.115 ;
        RECT 111.310 158.035 112.660 158.070 ;
      LAYER nwell ;
        RECT 71.060 154.935 119.740 157.765 ;
      LAYER pwell ;
        RECT 71.255 153.735 72.625 154.545 ;
        RECT 78.065 154.415 78.995 154.635 ;
        RECT 81.825 154.415 82.745 154.645 ;
        RECT 73.555 153.735 82.745 154.415 ;
        RECT 82.755 153.735 84.125 154.545 ;
        RECT 84.145 153.820 84.575 154.605 ;
        RECT 84.690 154.415 85.610 154.645 ;
        RECT 88.370 154.415 89.290 154.645 ;
        RECT 96.465 154.415 97.395 154.635 ;
        RECT 100.225 154.415 101.145 154.645 ;
        RECT 104.670 154.415 105.580 154.635 ;
        RECT 107.115 154.415 108.465 154.645 ;
        RECT 84.690 153.735 88.155 154.415 ;
        RECT 88.370 153.735 91.835 154.415 ;
        RECT 91.955 153.735 101.145 154.415 ;
        RECT 101.155 153.735 108.465 154.415 ;
        RECT 108.525 153.735 109.875 154.645 ;
        RECT 109.905 153.820 110.335 154.605 ;
        RECT 114.330 154.415 115.240 154.635 ;
        RECT 116.775 154.415 118.125 154.645 ;
        RECT 110.815 153.735 118.125 154.415 ;
        RECT 118.175 153.735 119.545 154.545 ;
      LAYER nwell ;
        RECT 17.405 152.860 22.575 153.700 ;
      LAYER pwell ;
        RECT 71.395 153.525 71.565 153.735 ;
        RECT 72.775 153.525 72.945 153.715 ;
        RECT 73.695 153.545 73.865 153.735 ;
        RECT 76.455 153.525 76.625 153.715 ;
        RECT 81.055 153.525 81.225 153.715 ;
        RECT 82.895 153.545 83.065 153.735 ;
        RECT 84.275 153.525 84.445 153.715 ;
        RECT 84.735 153.525 84.905 153.715 ;
        RECT 87.490 153.575 87.610 153.685 ;
        RECT 87.955 153.545 88.125 153.735 ;
        RECT 91.635 153.545 91.805 153.735 ;
        RECT 92.095 153.545 92.265 153.735 ;
        RECT 96.695 153.525 96.865 153.715 ;
        RECT 97.615 153.525 97.785 153.715 ;
        RECT 100.370 153.575 100.490 153.685 ;
        RECT 101.295 153.545 101.465 153.735 ;
        RECT 103.595 153.525 103.765 153.715 ;
        RECT 104.055 153.525 104.225 153.715 ;
        RECT 109.575 153.545 109.745 153.735 ;
        RECT 110.490 153.575 110.610 153.685 ;
        RECT 110.955 153.545 111.125 153.735 ;
        RECT 111.410 153.575 111.530 153.685 ;
        RECT 111.875 153.525 112.045 153.715 ;
        RECT 115.555 153.525 115.725 153.715 ;
        RECT 117.845 153.525 118.015 153.715 ;
        RECT 119.235 153.525 119.405 153.735 ;
      LAYER nwell ;
        RECT 17.410 150.285 22.530 152.860 ;
      LAYER pwell ;
        RECT 71.255 152.715 72.625 153.525 ;
        RECT 72.635 152.715 76.305 153.525 ;
        RECT 76.315 152.715 77.685 153.525 ;
        RECT 77.790 152.845 81.255 153.525 ;
        RECT 77.790 152.615 78.710 152.845 ;
        RECT 81.375 152.615 84.545 153.525 ;
        RECT 84.595 152.715 87.345 153.525 ;
        RECT 87.900 152.845 97.005 153.525 ;
        RECT 97.025 152.655 97.455 153.440 ;
        RECT 97.475 152.715 100.225 153.525 ;
        RECT 100.825 152.615 103.825 153.525 ;
        RECT 103.915 152.845 111.225 153.525 ;
        RECT 111.845 152.845 115.310 153.525 ;
        RECT 107.430 152.625 108.340 152.845 ;
        RECT 109.875 152.615 111.225 152.845 ;
        RECT 114.390 152.615 115.310 152.845 ;
        RECT 115.415 152.715 116.785 153.525 ;
        RECT 116.795 152.745 118.165 153.525 ;
        RECT 118.175 152.715 119.545 153.525 ;
      LAYER nwell ;
        RECT 71.060 149.495 119.740 152.325 ;
      LAYER pwell ;
        RECT 71.255 148.295 72.625 149.105 ;
        RECT 72.635 148.295 78.145 149.105 ;
        RECT 78.155 148.295 80.905 149.105 ;
        RECT 80.915 148.295 82.285 149.075 ;
        RECT 82.295 148.295 84.125 149.105 ;
        RECT 84.145 148.380 84.575 149.165 ;
        RECT 89.105 148.975 90.035 149.195 ;
        RECT 92.865 148.975 93.785 149.205 ;
        RECT 84.595 148.295 93.785 148.975 ;
        RECT 93.795 148.295 96.545 149.105 ;
        RECT 97.025 148.380 97.455 149.165 ;
        RECT 97.475 148.295 102.985 149.105 ;
        RECT 102.995 148.295 104.365 149.105 ;
        RECT 104.375 148.295 105.745 149.075 ;
        RECT 105.835 148.295 108.835 149.205 ;
        RECT 109.905 148.380 110.335 149.165 ;
        RECT 110.450 148.975 111.370 149.205 ;
        RECT 114.590 148.975 115.510 149.205 ;
        RECT 110.450 148.295 113.915 148.975 ;
        RECT 114.590 148.295 118.055 148.975 ;
        RECT 118.175 148.295 119.545 149.105 ;
        RECT 71.395 148.105 71.565 148.295 ;
        RECT 72.775 148.105 72.945 148.295 ;
        RECT 78.295 148.105 78.465 148.295 ;
        RECT 81.975 148.105 82.145 148.295 ;
        RECT 82.435 148.105 82.605 148.295 ;
        RECT 84.735 148.105 84.905 148.295 ;
        RECT 93.935 148.105 94.105 148.295 ;
        RECT 96.690 148.135 96.810 148.245 ;
        RECT 97.615 148.105 97.785 148.295 ;
        RECT 103.135 148.105 103.305 148.295 ;
        RECT 104.515 148.105 104.685 148.295 ;
        RECT 105.895 148.105 106.065 148.295 ;
        RECT 109.125 148.140 109.285 148.250 ;
        RECT 113.715 148.105 113.885 148.295 ;
        RECT 114.170 148.135 114.290 148.245 ;
        RECT 117.855 148.105 118.025 148.295 ;
        RECT 119.235 148.105 119.405 148.295 ;
      LAYER nwell ;
        RECT 14.250 136.535 31.270 137.965 ;
        RECT 14.250 133.205 15.680 136.535 ;
      LAYER pwell ;
        RECT 23.120 136.340 27.250 136.345 ;
        RECT 23.120 136.335 29.275 136.340 ;
        RECT 17.030 133.245 29.275 136.335 ;
        RECT 17.030 133.235 23.200 133.245 ;
        RECT 27.165 133.240 29.275 133.245 ;
      LAYER nwell ;
        RECT 29.760 133.205 31.270 136.535 ;
        RECT 14.250 131.775 31.270 133.205 ;
        RECT 17.185 114.890 22.355 115.730 ;
        RECT 17.190 112.315 22.310 114.890 ;
        RECT 14.030 98.565 31.050 99.995 ;
        RECT 14.030 95.235 15.460 98.565 ;
      LAYER pwell ;
        RECT 22.900 98.370 27.030 98.375 ;
        RECT 22.900 98.365 29.055 98.370 ;
        RECT 16.810 95.275 29.055 98.365 ;
        RECT 16.810 95.265 22.980 95.275 ;
        RECT 26.945 95.270 29.055 95.275 ;
      LAYER nwell ;
        RECT 29.540 95.235 31.050 98.565 ;
        RECT 14.030 93.805 31.050 95.235 ;
      LAYER pwell ;
        RECT 91.205 88.835 91.375 89.025 ;
        RECT 92.585 88.835 92.755 89.025 ;
        RECT 98.105 88.835 98.275 89.025 ;
        RECT 103.620 88.885 103.740 88.995 ;
        RECT 106.845 88.835 107.015 89.025 ;
        RECT 107.305 88.835 107.475 89.025 ;
        RECT 112.825 88.835 112.995 89.025 ;
        RECT 116.500 88.885 116.620 88.995 ;
        RECT 117.425 88.835 117.595 89.025 ;
        RECT 122.945 88.835 123.115 89.025 ;
        RECT 128.465 88.835 128.635 89.025 ;
        RECT 130.305 88.835 130.475 89.025 ;
        RECT 135.825 88.835 135.995 89.025 ;
        RECT 139.500 88.885 139.620 88.995 ;
        RECT 139.965 88.835 140.135 89.025 ;
        RECT 143.185 88.835 143.355 89.025 ;
        RECT 148.700 88.885 148.820 88.995 ;
        RECT 150.545 88.835 150.715 89.025 ;
        RECT 151.925 88.835 152.095 89.025 ;
        RECT 91.065 88.025 92.435 88.835 ;
        RECT 92.445 88.025 97.955 88.835 ;
        RECT 97.965 88.025 103.475 88.835 ;
        RECT 103.955 87.965 104.385 88.750 ;
        RECT 104.415 88.155 107.155 88.835 ;
        RECT 107.165 88.025 112.675 88.835 ;
        RECT 112.685 88.025 116.355 88.835 ;
        RECT 116.835 87.965 117.265 88.750 ;
        RECT 117.285 88.025 122.795 88.835 ;
        RECT 122.805 88.025 128.315 88.835 ;
        RECT 128.325 88.025 129.695 88.835 ;
        RECT 129.715 87.965 130.145 88.750 ;
        RECT 130.165 88.025 135.675 88.835 ;
        RECT 135.685 88.025 139.355 88.835 ;
        RECT 139.825 88.155 142.565 88.835 ;
        RECT 142.595 87.965 143.025 88.750 ;
        RECT 143.045 88.025 148.555 88.835 ;
        RECT 149.025 88.155 150.855 88.835 ;
        RECT 150.865 88.025 152.235 88.835 ;
      LAYER nwell ;
        RECT 90.870 84.805 152.430 87.635 ;
      LAYER pwell ;
        RECT 91.065 83.605 92.435 84.415 ;
        RECT 92.445 83.605 97.955 84.415 ;
        RECT 97.965 83.605 103.475 84.415 ;
        RECT 103.955 83.690 104.385 84.475 ;
        RECT 104.405 83.605 109.915 84.415 ;
        RECT 109.925 83.605 115.435 84.415 ;
        RECT 115.445 83.605 120.955 84.415 ;
        RECT 121.905 83.605 123.255 84.515 ;
        RECT 123.265 83.605 125.095 84.415 ;
        RECT 125.105 83.605 126.475 84.385 ;
        RECT 126.485 83.605 129.235 84.415 ;
        RECT 129.715 83.690 130.145 84.475 ;
        RECT 131.305 84.425 132.255 84.515 ;
        RECT 130.325 83.605 132.255 84.425 ;
        RECT 132.465 83.605 133.835 84.415 ;
        RECT 133.845 83.605 135.215 84.385 ;
        RECT 135.225 83.605 136.595 84.415 ;
        RECT 141.115 84.285 142.045 84.505 ;
        RECT 144.875 84.285 146.215 84.515 ;
        RECT 136.605 83.605 146.215 84.285 ;
        RECT 146.265 83.605 149.935 84.415 ;
        RECT 150.865 83.605 152.235 84.415 ;
        RECT 91.205 83.395 91.375 83.605 ;
        RECT 92.585 83.395 92.755 83.605 ;
        RECT 98.105 83.395 98.275 83.605 ;
        RECT 103.625 83.555 103.795 83.585 ;
        RECT 103.620 83.445 103.795 83.555 ;
        RECT 103.625 83.395 103.795 83.445 ;
        RECT 104.545 83.415 104.715 83.605 ;
        RECT 109.145 83.395 109.315 83.585 ;
        RECT 110.065 83.415 110.235 83.605 ;
        RECT 112.835 83.440 112.995 83.550 ;
        RECT 113.745 83.395 113.915 83.585 ;
        RECT 115.585 83.415 115.755 83.605 ;
        RECT 116.045 83.395 116.215 83.585 ;
        RECT 116.500 83.445 116.620 83.555 ;
        RECT 119.265 83.395 119.435 83.585 ;
        RECT 119.735 83.440 119.895 83.550 ;
        RECT 120.645 83.415 120.815 83.585 ;
        RECT 121.115 83.450 121.275 83.560 ;
        RECT 122.020 83.415 122.190 83.605 ;
        RECT 120.650 83.395 120.815 83.415 ;
        RECT 122.945 83.395 123.115 83.585 ;
        RECT 123.405 83.415 123.575 83.605 ;
        RECT 126.165 83.415 126.335 83.605 ;
        RECT 126.625 83.415 126.795 83.605 ;
        RECT 130.325 83.585 130.475 83.605 ;
        RECT 129.380 83.445 129.500 83.555 ;
        RECT 130.305 83.415 130.475 83.585 ;
        RECT 132.605 83.555 132.775 83.605 ;
        RECT 132.600 83.445 132.775 83.555 ;
        RECT 132.605 83.415 132.775 83.445 ;
        RECT 133.985 83.415 134.155 83.605 ;
        RECT 135.365 83.395 135.535 83.605 ;
        RECT 135.825 83.395 135.995 83.585 ;
        RECT 136.745 83.415 136.915 83.605 ;
        RECT 137.660 83.445 137.780 83.555 ;
        RECT 139.045 83.395 139.215 83.585 ;
        RECT 139.505 83.395 139.675 83.585 ;
        RECT 142.260 83.445 142.380 83.555 ;
        RECT 144.105 83.395 144.275 83.585 ;
        RECT 144.565 83.395 144.735 83.585 ;
        RECT 146.405 83.415 146.575 83.605 ;
        RECT 150.095 83.440 150.255 83.560 ;
        RECT 151.925 83.395 152.095 83.605 ;
        RECT 91.065 82.585 92.435 83.395 ;
        RECT 92.445 82.585 97.955 83.395 ;
        RECT 97.965 82.585 103.475 83.395 ;
        RECT 103.485 82.585 108.995 83.395 ;
        RECT 109.005 82.585 112.675 83.395 ;
        RECT 113.615 82.485 114.965 83.395 ;
        RECT 114.985 82.615 116.355 83.395 ;
        RECT 116.835 82.525 117.265 83.310 ;
        RECT 117.285 82.715 119.575 83.395 ;
        RECT 120.650 82.715 122.485 83.395 ;
        RECT 122.805 82.715 132.415 83.395 ;
        RECT 117.285 82.485 118.205 82.715 ;
        RECT 121.555 82.485 122.485 82.715 ;
        RECT 127.315 82.495 128.245 82.715 ;
        RECT 131.075 82.485 132.415 82.715 ;
        RECT 132.925 82.485 135.675 83.395 ;
        RECT 135.685 82.585 137.515 83.395 ;
        RECT 137.995 82.485 139.345 83.395 ;
        RECT 139.365 82.585 142.115 83.395 ;
        RECT 142.595 82.525 143.025 83.310 ;
        RECT 143.055 82.485 144.405 83.395 ;
        RECT 144.425 82.585 149.935 83.395 ;
        RECT 150.865 82.585 152.235 83.395 ;
      LAYER nwell ;
        RECT 90.870 79.365 152.430 82.195 ;
      LAYER pwell ;
        RECT 91.065 78.165 92.435 78.975 ;
        RECT 92.445 78.165 97.955 78.975 ;
        RECT 97.965 78.165 103.475 78.975 ;
        RECT 103.955 78.250 104.385 79.035 ;
        RECT 104.405 78.165 109.915 78.975 ;
        RECT 115.355 78.845 116.285 79.065 ;
        RECT 119.115 78.845 120.455 79.075 ;
        RECT 122.795 78.845 123.715 79.075 ;
        RECT 110.845 78.165 120.455 78.845 ;
        RECT 121.425 78.165 123.715 78.845 ;
        RECT 124.745 78.165 127.855 79.075 ;
        RECT 127.875 78.165 129.225 79.075 ;
        RECT 129.715 78.250 130.145 79.035 ;
        RECT 131.085 78.165 134.295 79.075 ;
        RECT 134.305 78.165 137.515 79.075 ;
        RECT 137.525 78.165 143.035 78.975 ;
        RECT 143.045 78.875 143.990 79.075 ;
        RECT 143.045 78.195 145.795 78.875 ;
        RECT 143.045 78.165 143.990 78.195 ;
        RECT 91.205 77.955 91.375 78.165 ;
        RECT 92.585 77.955 92.755 78.165 ;
        RECT 98.105 77.955 98.275 78.165 ;
        RECT 103.625 78.115 103.795 78.145 ;
        RECT 103.620 78.005 103.795 78.115 ;
        RECT 103.625 77.955 103.795 78.005 ;
        RECT 104.545 77.975 104.715 78.165 ;
        RECT 107.305 77.955 107.475 78.145 ;
        RECT 109.605 77.955 109.775 78.145 ;
        RECT 110.065 77.955 110.235 78.145 ;
        RECT 110.985 77.975 111.155 78.165 ;
        RECT 115.585 77.955 115.755 78.145 ;
        RECT 117.425 77.955 117.595 78.145 ;
        RECT 118.805 77.955 118.975 78.145 ;
        RECT 120.655 78.010 120.815 78.120 ;
        RECT 121.565 77.975 121.735 78.165 ;
        RECT 122.025 77.955 122.195 78.145 ;
        RECT 122.485 77.955 122.655 78.145 ;
        RECT 123.875 78.010 124.035 78.120 ;
        RECT 124.785 77.975 124.955 78.165 ;
        RECT 128.005 77.955 128.175 78.165 ;
        RECT 129.380 78.005 129.500 78.115 ;
        RECT 130.315 78.010 130.475 78.120 ;
        RECT 131.225 77.975 131.395 78.165 ;
        RECT 134.435 78.145 134.605 78.165 ;
        RECT 134.435 77.975 134.615 78.145 ;
        RECT 134.445 77.955 134.615 77.975 ;
        RECT 134.905 77.955 135.075 78.145 ;
        RECT 137.665 77.975 137.835 78.165 ;
        RECT 138.125 77.955 138.295 78.145 ;
        RECT 140.890 77.955 141.060 78.145 ;
        RECT 143.185 77.955 143.355 78.145 ;
        RECT 145.480 77.975 145.650 78.195 ;
        RECT 145.805 78.165 149.475 78.975 ;
        RECT 149.485 78.165 150.855 78.975 ;
        RECT 150.865 78.165 152.235 78.975 ;
        RECT 145.945 77.975 146.115 78.165 ;
        RECT 146.405 77.955 146.575 78.145 ;
        RECT 147.785 77.955 147.955 78.145 ;
        RECT 149.625 77.975 149.795 78.165 ;
        RECT 150.540 78.005 150.660 78.115 ;
        RECT 151.925 77.955 152.095 78.165 ;
        RECT 91.065 77.145 92.435 77.955 ;
        RECT 92.445 77.145 97.955 77.955 ;
        RECT 97.965 77.145 103.475 77.955 ;
        RECT 103.485 77.145 107.155 77.955 ;
        RECT 107.165 77.145 108.535 77.955 ;
        RECT 108.545 77.175 109.915 77.955 ;
        RECT 109.925 77.145 115.435 77.955 ;
        RECT 115.445 77.145 116.815 77.955 ;
        RECT 116.835 77.085 117.265 77.870 ;
        RECT 117.285 77.145 118.655 77.955 ;
        RECT 118.665 77.275 120.955 77.955 ;
        RECT 120.035 77.045 120.955 77.275 ;
        RECT 120.975 77.045 122.325 77.955 ;
        RECT 122.345 77.145 127.855 77.955 ;
        RECT 127.865 77.145 131.535 77.955 ;
        RECT 131.545 77.275 134.755 77.955 ;
        RECT 131.545 77.045 132.680 77.275 ;
        RECT 134.765 77.045 137.975 77.955 ;
        RECT 137.985 77.145 140.735 77.955 ;
        RECT 140.745 77.045 142.575 77.955 ;
        RECT 142.595 77.085 143.025 77.870 ;
        RECT 143.145 77.045 146.255 77.955 ;
        RECT 146.275 77.045 147.625 77.955 ;
        RECT 147.645 77.145 150.395 77.955 ;
        RECT 150.865 77.145 152.235 77.955 ;
      LAYER nwell ;
        RECT 90.870 73.925 152.430 76.755 ;
      LAYER pwell ;
        RECT 91.065 72.725 92.435 73.535 ;
        RECT 92.445 72.725 97.955 73.535 ;
        RECT 97.965 72.725 103.475 73.535 ;
        RECT 103.955 72.810 104.385 73.595 ;
        RECT 108.915 73.405 109.845 73.625 ;
        RECT 112.565 73.405 114.775 73.635 ;
        RECT 104.405 72.725 114.775 73.405 ;
        RECT 115.085 72.725 118.195 73.635 ;
        RECT 118.205 72.725 119.575 73.535 ;
        RECT 119.585 72.725 122.505 73.635 ;
        RECT 122.805 72.725 125.555 73.535 ;
        RECT 126.335 73.405 127.265 73.635 ;
        RECT 126.335 72.725 128.170 73.405 ;
        RECT 128.325 72.725 129.695 73.535 ;
        RECT 129.715 72.810 130.145 73.595 ;
        RECT 130.625 72.725 133.835 73.635 ;
        RECT 133.845 72.725 139.355 73.535 ;
        RECT 139.365 72.725 140.735 73.535 ;
        RECT 140.755 72.725 142.105 73.635 ;
        RECT 142.605 72.725 143.955 73.635 ;
        RECT 143.965 72.725 147.440 73.635 ;
        RECT 147.645 72.725 150.395 73.535 ;
        RECT 150.865 72.725 152.235 73.535 ;
        RECT 91.205 72.515 91.375 72.725 ;
        RECT 92.585 72.515 92.755 72.725 ;
        RECT 98.105 72.515 98.275 72.725 ;
        RECT 103.625 72.675 103.795 72.705 ;
        RECT 103.620 72.565 103.795 72.675 ;
        RECT 103.625 72.515 103.795 72.565 ;
        RECT 104.545 72.535 104.715 72.725 ;
        RECT 107.305 72.515 107.475 72.705 ;
        RECT 108.685 72.515 108.855 72.705 ;
        RECT 110.065 72.515 110.235 72.705 ;
        RECT 113.745 72.515 113.915 72.705 ;
        RECT 115.125 72.515 115.295 72.725 ;
        RECT 118.345 72.535 118.515 72.725 ;
        RECT 119.730 72.705 119.900 72.725 ;
        RECT 119.725 72.535 119.900 72.705 ;
        RECT 119.725 72.515 119.895 72.535 ;
        RECT 120.185 72.515 120.355 72.705 ;
        RECT 121.565 72.515 121.735 72.705 ;
        RECT 122.945 72.535 123.115 72.725 ;
        RECT 128.005 72.705 128.170 72.725 ;
        RECT 125.700 72.565 125.820 72.675 ;
        RECT 126.160 72.515 126.330 72.705 ;
        RECT 126.625 72.515 126.795 72.705 ;
        RECT 128.005 72.535 128.175 72.705 ;
        RECT 128.465 72.515 128.635 72.725 ;
        RECT 130.300 72.565 130.420 72.675 ;
        RECT 130.755 72.535 130.925 72.725 ;
        RECT 132.145 72.515 132.315 72.705 ;
        RECT 133.525 72.515 133.695 72.705 ;
        RECT 133.985 72.535 134.155 72.725 ;
        RECT 137.665 72.515 137.835 72.705 ;
        RECT 138.120 72.565 138.240 72.675 ;
        RECT 139.505 72.515 139.675 72.725 ;
        RECT 139.965 72.515 140.135 72.705 ;
        RECT 141.805 72.535 141.975 72.725 ;
        RECT 142.260 72.565 142.380 72.675 ;
        RECT 142.720 72.535 142.890 72.725 ;
        RECT 91.065 71.705 92.435 72.515 ;
        RECT 92.445 71.705 97.955 72.515 ;
        RECT 97.965 71.705 103.475 72.515 ;
        RECT 103.485 71.705 107.155 72.515 ;
        RECT 107.165 71.705 108.535 72.515 ;
        RECT 108.555 71.605 109.905 72.515 ;
        RECT 109.925 71.705 113.595 72.515 ;
        RECT 113.605 71.705 114.975 72.515 ;
        RECT 115.000 71.605 116.815 72.515 ;
        RECT 116.835 71.645 117.265 72.430 ;
        RECT 117.285 71.835 120.035 72.515 ;
        RECT 117.285 71.605 118.215 71.835 ;
        RECT 120.045 71.705 121.415 72.515 ;
        RECT 121.535 71.835 125.000 72.515 ;
        RECT 124.080 71.605 125.000 71.835 ;
        RECT 125.125 71.605 126.475 72.515 ;
        RECT 126.500 71.605 128.315 72.515 ;
        RECT 128.325 71.705 131.995 72.515 ;
        RECT 132.005 71.705 133.375 72.515 ;
        RECT 133.465 71.605 136.465 72.515 ;
        RECT 136.615 71.605 137.965 72.515 ;
        RECT 138.455 71.605 139.805 72.515 ;
        RECT 139.825 71.835 142.575 72.515 ;
        RECT 143.190 72.485 143.360 72.705 ;
        RECT 144.110 72.535 144.280 72.725 ;
        RECT 147.785 72.535 147.955 72.725 ;
        RECT 150.570 72.675 150.740 72.705 ;
        RECT 150.540 72.565 150.740 72.675 ;
        RECT 150.570 72.535 150.740 72.565 ;
        RECT 150.570 72.515 150.680 72.535 ;
        RECT 151.925 72.515 152.095 72.725 ;
        RECT 145.320 72.485 146.255 72.515 ;
        RECT 141.645 71.605 142.575 71.835 ;
        RECT 142.595 71.645 143.025 72.430 ;
        RECT 143.190 72.285 146.255 72.485 ;
        RECT 143.045 71.805 146.255 72.285 ;
        RECT 143.045 71.605 143.975 71.805 ;
        RECT 145.305 71.605 146.255 71.805 ;
        RECT 146.265 71.835 150.680 72.515 ;
        RECT 146.265 71.605 150.195 71.835 ;
        RECT 150.865 71.705 152.235 72.515 ;
      LAYER nwell ;
        RECT 21.650 68.590 22.740 68.990 ;
        RECT 24.070 68.590 25.600 68.990 ;
        RECT 29.400 68.590 30.930 68.990 ;
        RECT 20.760 68.580 26.360 68.590 ;
        RECT 28.630 68.580 31.690 68.590 ;
        RECT 33.650 68.580 34.495 68.585 ;
        RECT 20.760 66.600 34.495 68.580 ;
        RECT 90.870 68.485 152.430 71.315 ;
      LAYER pwell ;
        RECT 91.065 67.285 92.435 68.095 ;
        RECT 92.445 67.285 97.955 68.095 ;
        RECT 97.965 67.285 100.715 68.095 ;
        RECT 101.185 67.285 102.555 68.065 ;
        RECT 102.565 67.285 103.935 68.095 ;
        RECT 103.955 67.370 104.385 68.155 ;
        RECT 104.405 67.285 109.915 68.095 ;
        RECT 115.355 67.965 116.285 68.185 ;
        RECT 119.115 67.965 120.455 68.195 ;
        RECT 110.845 67.285 120.455 67.965 ;
        RECT 120.705 68.105 121.655 68.195 ;
        RECT 120.705 67.285 122.635 68.105 ;
        RECT 122.805 67.285 128.315 68.095 ;
        RECT 128.325 67.285 129.695 68.095 ;
        RECT 129.715 67.370 130.145 68.155 ;
        RECT 130.165 67.285 131.995 68.095 ;
        RECT 133.825 67.965 134.755 68.195 ;
        RECT 136.570 67.995 137.515 68.195 ;
        RECT 139.330 67.995 140.275 68.195 ;
        RECT 132.005 67.285 134.755 67.965 ;
        RECT 134.765 67.315 137.515 67.995 ;
        RECT 137.525 67.315 140.275 67.995 ;
        RECT 91.205 67.075 91.375 67.285 ;
        RECT 92.585 67.075 92.755 67.285 ;
        RECT 98.105 67.235 98.275 67.285 ;
        RECT 98.100 67.125 98.275 67.235 ;
        RECT 98.105 67.095 98.275 67.125 ;
        RECT 98.565 67.075 98.735 67.265 ;
        RECT 100.860 67.125 100.980 67.235 ;
        RECT 102.245 67.095 102.415 67.285 ;
        RECT 102.705 67.095 102.875 67.285 ;
        RECT 104.545 67.095 104.715 67.285 ;
        RECT 109.145 67.075 109.315 67.265 ;
        RECT 109.605 67.075 109.775 67.265 ;
        RECT 110.075 67.130 110.235 67.240 ;
        RECT 110.985 67.095 111.155 67.285 ;
        RECT 122.485 67.265 122.635 67.285 ;
        RECT 115.125 67.075 115.295 67.265 ;
        RECT 116.500 67.125 116.620 67.235 ;
        RECT 117.425 67.075 117.595 67.265 ;
        RECT 121.115 67.120 121.275 67.230 ;
        RECT 122.485 67.095 122.655 67.265 ;
        RECT 122.945 67.075 123.115 67.285 ;
        RECT 123.415 67.120 123.575 67.230 ;
        RECT 124.325 67.075 124.495 67.265 ;
        RECT 128.465 67.095 128.635 67.285 ;
        RECT 130.305 67.095 130.475 67.285 ;
        RECT 132.145 67.095 132.315 67.285 ;
        RECT 133.520 67.125 133.640 67.235 ;
        RECT 133.990 67.075 134.160 67.265 ;
        RECT 134.910 67.095 135.080 67.315 ;
        RECT 136.570 67.285 137.515 67.315 ;
        RECT 135.825 67.075 135.995 67.265 ;
        RECT 137.670 67.235 137.840 67.315 ;
        RECT 139.330 67.285 140.275 67.315 ;
        RECT 140.285 67.285 142.115 68.095 ;
        RECT 142.585 67.285 146.240 68.195 ;
        RECT 146.265 67.995 147.210 68.195 ;
        RECT 146.265 67.315 149.015 67.995 ;
        RECT 146.265 67.285 147.210 67.315 ;
        RECT 137.660 67.125 137.840 67.235 ;
        RECT 137.670 67.095 137.840 67.125 ;
        RECT 138.125 67.075 138.295 67.265 ;
        RECT 140.425 67.095 140.595 67.285 ;
        RECT 142.260 67.125 142.380 67.235 ;
        RECT 142.730 67.095 142.900 67.285 ;
      LAYER nwell ;
        RECT 20.760 65.125 33.995 66.600 ;
      LAYER pwell ;
        RECT 91.065 66.265 92.435 67.075 ;
        RECT 92.445 66.265 97.955 67.075 ;
        RECT 98.425 66.395 108.035 67.075 ;
        RECT 102.935 66.175 103.865 66.395 ;
        RECT 106.695 66.165 108.035 66.395 ;
        RECT 108.095 66.165 109.445 67.075 ;
        RECT 109.465 66.265 114.975 67.075 ;
        RECT 114.995 66.165 116.345 67.075 ;
        RECT 116.835 66.205 117.265 66.990 ;
        RECT 117.285 66.265 120.955 67.075 ;
        RECT 121.895 66.165 123.245 67.075 ;
        RECT 124.185 66.395 133.375 67.075 ;
        RECT 128.695 66.175 129.625 66.395 ;
        RECT 132.455 66.165 133.375 66.395 ;
        RECT 133.845 66.165 135.675 67.075 ;
        RECT 135.685 66.265 137.515 67.075 ;
        RECT 137.985 66.165 142.045 67.075 ;
        RECT 143.050 67.045 144.450 67.075 ;
        RECT 145.940 67.045 146.110 67.265 ;
        RECT 146.405 67.075 146.575 67.265 ;
        RECT 148.700 67.095 148.870 67.315 ;
        RECT 149.025 67.285 150.855 68.095 ;
        RECT 150.865 67.285 152.235 68.095 ;
        RECT 149.165 67.095 149.335 67.285 ;
        RECT 150.095 67.120 150.255 67.230 ;
        RECT 151.925 67.075 152.095 67.285 ;
        RECT 142.595 66.205 143.025 66.990 ;
        RECT 143.050 66.365 146.255 67.045 ;
        RECT 143.050 66.165 144.450 66.365 ;
        RECT 146.265 66.265 149.935 67.075 ;
        RECT 150.865 66.265 152.235 67.075 ;
      LAYER nwell ;
        RECT 21.660 65.080 33.995 65.125 ;
        RECT 23.295 65.045 33.995 65.080 ;
        RECT 23.300 65.040 33.995 65.045 ;
        RECT 31.855 64.980 33.995 65.040 ;
        RECT 90.870 63.045 152.430 65.875 ;
      LAYER pwell ;
        RECT 91.065 61.845 92.435 62.655 ;
        RECT 92.485 62.525 93.825 62.755 ;
        RECT 96.655 62.525 97.585 62.745 ;
        RECT 92.485 61.845 102.095 62.525 ;
        RECT 102.115 61.845 103.465 62.755 ;
        RECT 103.955 61.930 104.385 62.715 ;
        RECT 104.405 61.845 105.775 62.655 ;
        RECT 105.785 62.525 106.715 62.755 ;
        RECT 109.465 62.525 110.395 62.755 ;
        RECT 117.195 62.525 118.125 62.745 ;
        RECT 120.955 62.525 121.875 62.755 ;
        RECT 105.785 61.845 109.455 62.525 ;
        RECT 109.465 61.845 112.215 62.525 ;
        RECT 112.685 61.845 121.875 62.525 ;
        RECT 121.980 62.525 122.900 62.755 ;
        RECT 121.980 61.845 125.445 62.525 ;
        RECT 126.495 61.845 127.845 62.755 ;
        RECT 127.865 61.845 129.695 62.655 ;
        RECT 129.715 61.930 130.145 62.715 ;
        RECT 130.165 61.845 135.675 62.655 ;
        RECT 135.685 61.845 141.195 62.655 ;
        RECT 142.125 61.845 143.475 62.755 ;
        RECT 143.505 61.845 146.255 62.655 ;
        RECT 146.275 61.845 147.625 62.755 ;
        RECT 147.645 61.845 150.395 62.655 ;
        RECT 150.865 61.845 152.235 62.655 ;
        RECT 91.205 61.635 91.375 61.845 ;
        RECT 101.785 61.825 101.955 61.845 ;
        RECT 92.585 61.635 92.755 61.825 ;
        RECT 96.275 61.680 96.435 61.790 ;
        RECT 97.180 61.635 97.350 61.825 ;
        RECT 101.780 61.655 101.955 61.825 ;
        RECT 103.165 61.655 103.335 61.845 ;
        RECT 103.620 61.685 103.740 61.795 ;
        RECT 104.545 61.655 104.715 61.845 ;
        RECT 101.780 61.635 101.950 61.655 ;
        RECT 91.065 60.825 92.435 61.635 ;
        RECT 92.445 60.825 96.115 61.635 ;
        RECT 97.065 60.725 98.415 61.635 ;
        RECT 98.620 60.725 102.095 61.635 ;
        RECT 102.105 61.605 103.040 61.635 ;
        RECT 105.000 61.605 105.170 61.825 ;
        RECT 105.465 61.635 105.635 61.825 ;
        RECT 108.225 61.635 108.395 61.825 ;
        RECT 109.145 61.655 109.315 61.845 ;
        RECT 111.905 61.655 112.075 61.845 ;
        RECT 112.360 61.685 112.480 61.795 ;
        RECT 112.825 61.655 112.995 61.845 ;
        RECT 113.740 61.685 113.860 61.795 ;
        RECT 114.205 61.635 114.375 61.825 ;
        RECT 117.425 61.635 117.595 61.825 ;
        RECT 125.245 61.655 125.415 61.845 ;
        RECT 125.715 61.690 125.875 61.800 ;
        RECT 126.625 61.635 126.795 61.845 ;
        RECT 128.005 61.655 128.175 61.845 ;
        RECT 130.305 61.655 130.475 61.845 ;
        RECT 132.145 61.635 132.315 61.825 ;
        RECT 135.825 61.655 135.995 61.845 ;
        RECT 137.665 61.635 137.835 61.825 ;
        RECT 141.345 61.635 141.515 61.825 ;
        RECT 142.270 61.655 142.440 61.845 ;
        RECT 143.185 61.635 143.355 61.825 ;
        RECT 143.645 61.655 143.815 61.845 ;
        RECT 145.945 61.635 146.115 61.825 ;
        RECT 147.325 61.655 147.495 61.845 ;
        RECT 147.785 61.655 147.955 61.845 ;
        RECT 150.545 61.795 150.715 61.825 ;
        RECT 150.540 61.685 150.715 61.795 ;
        RECT 150.545 61.635 150.715 61.685 ;
        RECT 151.925 61.635 152.095 61.845 ;
        RECT 102.105 61.405 105.170 61.605 ;
        RECT 102.105 60.925 105.315 61.405 ;
        RECT 102.105 60.725 103.055 60.925 ;
        RECT 104.385 60.725 105.315 60.925 ;
        RECT 105.335 60.725 108.065 61.635 ;
        RECT 108.085 60.825 113.595 61.635 ;
        RECT 114.075 60.725 116.805 61.635 ;
        RECT 116.835 60.765 117.265 61.550 ;
        RECT 117.285 60.955 126.390 61.635 ;
        RECT 126.485 60.825 131.995 61.635 ;
        RECT 132.005 60.825 137.515 61.635 ;
        RECT 137.525 60.825 141.195 61.635 ;
        RECT 141.205 60.825 142.575 61.635 ;
        RECT 142.595 60.765 143.025 61.550 ;
        RECT 143.045 60.825 145.795 61.635 ;
        RECT 145.815 60.725 147.165 61.635 ;
        RECT 147.280 60.955 150.745 61.635 ;
        RECT 147.280 60.725 148.200 60.955 ;
        RECT 150.865 60.825 152.235 61.635 ;
      LAYER nwell ;
        RECT 90.870 57.605 152.430 60.435 ;
      LAYER pwell ;
        RECT 91.065 56.405 92.435 57.215 ;
        RECT 92.445 56.405 96.115 57.215 ;
        RECT 96.585 56.405 98.415 57.315 ;
        RECT 98.625 57.225 99.575 57.315 ;
        RECT 100.925 57.225 101.875 57.315 ;
        RECT 98.625 56.405 100.555 57.225 ;
        RECT 100.925 56.405 102.855 57.225 ;
        RECT 103.955 56.490 104.385 57.275 ;
        RECT 104.405 56.405 109.915 57.215 ;
        RECT 109.925 56.405 111.755 57.215 ;
        RECT 111.850 56.405 120.955 57.085 ;
        RECT 120.965 56.405 124.635 57.215 ;
        RECT 125.115 56.405 126.465 57.315 ;
        RECT 126.485 56.405 127.855 57.185 ;
        RECT 127.865 56.405 129.695 57.215 ;
        RECT 129.715 56.490 130.145 57.275 ;
        RECT 131.215 57.085 132.145 57.315 ;
        RECT 130.310 56.405 132.145 57.085 ;
        RECT 132.925 56.405 134.295 57.185 ;
        RECT 134.305 56.405 139.815 57.215 ;
        RECT 139.825 56.405 141.195 57.215 ;
        RECT 145.715 57.085 146.645 57.305 ;
        RECT 149.475 57.085 150.395 57.315 ;
        RECT 141.205 56.405 150.395 57.085 ;
        RECT 150.865 56.405 152.235 57.215 ;
        RECT 91.205 56.195 91.375 56.405 ;
        RECT 92.585 56.195 92.755 56.405 ;
        RECT 96.260 56.245 96.380 56.355 ;
        RECT 98.100 56.215 98.270 56.405 ;
        RECT 100.405 56.385 100.555 56.405 ;
        RECT 102.705 56.385 102.855 56.405 ;
        RECT 98.570 56.195 98.740 56.385 ;
        RECT 99.945 56.195 100.115 56.385 ;
        RECT 100.405 56.215 100.575 56.385 ;
        RECT 102.705 56.215 102.875 56.385 ;
        RECT 103.175 56.250 103.335 56.360 ;
        RECT 104.545 56.215 104.715 56.405 ;
        RECT 105.465 56.195 105.635 56.385 ;
        RECT 110.065 56.215 110.235 56.405 ;
        RECT 110.985 56.195 111.155 56.385 ;
        RECT 91.065 55.385 92.435 56.195 ;
        RECT 92.445 55.385 97.955 56.195 ;
        RECT 98.425 55.285 99.775 56.195 ;
        RECT 99.805 55.385 105.315 56.195 ;
        RECT 105.325 55.385 110.835 56.195 ;
        RECT 110.845 55.385 112.215 56.195 ;
        RECT 112.370 56.165 112.540 56.385 ;
        RECT 116.505 56.195 116.675 56.385 ;
        RECT 117.435 56.240 117.595 56.350 ;
        RECT 118.345 56.195 118.515 56.385 ;
        RECT 119.725 56.195 119.895 56.385 ;
        RECT 120.645 56.215 120.815 56.405 ;
        RECT 121.105 56.215 121.275 56.405 ;
        RECT 124.780 56.245 124.900 56.355 ;
        RECT 126.165 56.215 126.335 56.405 ;
        RECT 126.625 56.215 126.795 56.405 ;
        RECT 128.005 56.215 128.175 56.405 ;
        RECT 130.310 56.385 130.475 56.405 ;
        RECT 130.305 56.215 130.475 56.385 ;
        RECT 130.765 56.195 130.935 56.385 ;
        RECT 131.220 56.245 131.340 56.355 ;
        RECT 131.685 56.195 131.855 56.385 ;
        RECT 132.600 56.245 132.720 56.355 ;
        RECT 133.985 56.215 134.155 56.405 ;
        RECT 134.445 56.215 134.615 56.405 ;
        RECT 139.965 56.215 140.135 56.405 ;
        RECT 141.345 56.215 141.515 56.405 ;
        RECT 141.805 56.195 141.975 56.385 ;
        RECT 142.260 56.245 142.380 56.355 ;
        RECT 143.185 56.195 143.355 56.385 ;
        RECT 145.940 56.245 146.060 56.355 ;
        RECT 146.405 56.195 146.575 56.385 ;
        RECT 147.785 56.195 147.955 56.385 ;
        RECT 150.540 56.245 150.660 56.355 ;
        RECT 151.925 56.195 152.095 56.405 ;
        RECT 114.500 56.165 115.435 56.195 ;
        RECT 112.370 55.965 115.435 56.165 ;
        RECT 112.225 55.485 115.435 55.965 ;
        RECT 112.225 55.285 113.155 55.485 ;
        RECT 114.485 55.285 115.435 55.485 ;
        RECT 115.445 55.415 116.815 56.195 ;
        RECT 116.835 55.325 117.265 56.110 ;
        RECT 118.215 55.285 119.565 56.195 ;
        RECT 119.585 55.385 121.415 56.195 ;
        RECT 121.465 55.515 131.075 56.195 ;
        RECT 131.545 55.515 140.735 56.195 ;
        RECT 121.465 55.285 122.805 55.515 ;
        RECT 125.635 55.295 126.565 55.515 ;
        RECT 136.055 55.295 136.985 55.515 ;
        RECT 139.815 55.285 140.735 55.515 ;
        RECT 140.755 55.285 142.105 56.195 ;
        RECT 142.595 55.325 143.025 56.110 ;
        RECT 143.045 55.385 145.795 56.195 ;
        RECT 146.275 55.285 147.625 56.195 ;
        RECT 147.645 55.385 150.395 56.195 ;
        RECT 150.865 55.385 152.235 56.195 ;
      LAYER nwell ;
        RECT 90.870 52.165 152.430 54.995 ;
      LAYER pwell ;
        RECT 91.065 50.965 92.435 51.775 ;
        RECT 96.955 51.645 97.885 51.865 ;
        RECT 100.715 51.645 101.635 51.875 ;
        RECT 92.445 50.965 101.635 51.645 ;
        RECT 101.655 50.965 103.005 51.875 ;
        RECT 103.955 51.050 104.385 51.835 ;
        RECT 104.405 50.965 106.235 51.775 ;
        RECT 107.295 51.645 108.225 51.875 ;
        RECT 106.390 50.965 108.225 51.645 ;
        RECT 109.005 50.965 110.375 51.745 ;
        RECT 111.895 51.645 112.825 51.875 ;
        RECT 117.655 51.645 118.585 51.865 ;
        RECT 121.415 51.645 122.335 51.875 ;
        RECT 124.405 51.785 125.355 51.875 ;
        RECT 110.990 50.965 112.825 51.645 ;
        RECT 113.145 50.965 122.335 51.645 ;
        RECT 123.425 50.965 125.355 51.785 ;
        RECT 125.565 51.675 126.495 51.875 ;
        RECT 127.825 51.675 128.775 51.875 ;
        RECT 125.565 51.195 128.775 51.675 ;
        RECT 125.710 50.995 128.775 51.195 ;
        RECT 129.715 51.050 130.145 51.835 ;
        RECT 131.085 51.675 132.035 51.875 ;
        RECT 133.365 51.675 134.295 51.875 ;
        RECT 131.085 51.195 134.295 51.675 ;
        RECT 134.305 51.645 135.225 51.875 ;
        RECT 136.605 51.675 137.535 51.875 ;
        RECT 138.865 51.675 139.815 51.875 ;
        RECT 91.205 50.755 91.375 50.965 ;
        RECT 92.585 50.755 92.755 50.965 ;
        RECT 96.265 50.755 96.435 50.945 ;
        RECT 98.565 50.755 98.735 50.945 ;
        RECT 99.945 50.755 100.115 50.945 ;
        RECT 100.405 50.755 100.575 50.945 ;
        RECT 102.245 50.775 102.415 50.945 ;
        RECT 102.705 50.775 102.875 50.965 ;
        RECT 103.175 50.810 103.335 50.920 ;
        RECT 104.545 50.915 104.715 50.965 ;
        RECT 106.390 50.945 106.555 50.965 ;
        RECT 104.540 50.805 104.715 50.915 ;
        RECT 104.545 50.775 104.715 50.805 ;
        RECT 106.385 50.775 106.555 50.945 ;
        RECT 102.265 50.755 102.415 50.775 ;
        RECT 106.845 50.755 107.015 50.945 ;
        RECT 107.305 50.755 107.475 50.945 ;
        RECT 108.680 50.805 108.800 50.915 ;
        RECT 110.065 50.775 110.235 50.965 ;
        RECT 110.990 50.945 111.155 50.965 ;
        RECT 110.520 50.805 110.640 50.915 ;
        RECT 110.985 50.775 111.155 50.945 ;
        RECT 113.285 50.775 113.455 50.965 ;
        RECT 123.425 50.945 123.575 50.965 ;
        RECT 117.425 50.755 117.595 50.945 ;
        RECT 122.495 50.810 122.655 50.920 ;
        RECT 122.945 50.755 123.115 50.945 ;
        RECT 123.405 50.775 123.575 50.945 ;
        RECT 125.710 50.775 125.880 50.995 ;
        RECT 127.840 50.965 128.775 50.995 ;
        RECT 131.085 50.995 134.150 51.195 ;
        RECT 131.085 50.965 132.020 50.995 ;
        RECT 126.625 50.775 126.795 50.945 ;
        RECT 126.630 50.755 126.795 50.775 ;
        RECT 128.925 50.755 129.095 50.945 ;
        RECT 130.315 50.810 130.475 50.920 ;
        RECT 131.680 50.805 131.800 50.915 ;
        RECT 132.145 50.755 132.315 50.945 ;
        RECT 133.980 50.775 134.150 50.995 ;
        RECT 134.305 50.965 136.595 51.645 ;
        RECT 136.605 51.195 139.815 51.675 ;
        RECT 136.750 50.995 139.815 51.195 ;
        RECT 135.365 50.775 135.535 50.945 ;
        RECT 136.285 50.775 136.455 50.965 ;
        RECT 136.750 50.775 136.920 50.995 ;
        RECT 138.880 50.965 139.815 50.995 ;
        RECT 139.825 50.965 141.195 51.745 ;
        RECT 145.715 51.645 146.645 51.865 ;
        RECT 149.475 51.645 150.395 51.875 ;
        RECT 141.205 50.965 150.395 51.645 ;
        RECT 150.865 50.965 152.235 51.775 ;
        RECT 135.370 50.755 135.535 50.775 ;
        RECT 137.665 50.755 137.835 50.945 ;
        RECT 139.965 50.775 140.135 50.965 ;
        RECT 141.345 50.755 141.515 50.965 ;
        RECT 143.185 50.755 143.355 50.945 ;
        RECT 150.570 50.915 150.740 50.945 ;
        RECT 145.940 50.805 146.060 50.915 ;
        RECT 150.540 50.805 150.740 50.915 ;
        RECT 150.570 50.775 150.740 50.805 ;
        RECT 150.570 50.755 150.680 50.775 ;
        RECT 151.925 50.755 152.095 50.965 ;
        RECT 91.065 49.945 92.435 50.755 ;
        RECT 92.445 49.945 96.115 50.755 ;
        RECT 96.125 49.945 97.495 50.755 ;
        RECT 97.505 49.975 98.875 50.755 ;
        RECT 98.895 49.845 100.245 50.755 ;
        RECT 100.265 49.945 102.095 50.755 ;
        RECT 102.265 49.935 104.195 50.755 ;
        RECT 103.245 49.845 104.195 49.935 ;
        RECT 104.865 50.075 107.155 50.755 ;
        RECT 107.165 50.075 116.775 50.755 ;
        RECT 104.865 49.845 105.785 50.075 ;
        RECT 111.675 49.855 112.605 50.075 ;
        RECT 115.435 49.845 116.775 50.075 ;
        RECT 116.835 49.885 117.265 50.670 ;
        RECT 117.285 49.945 122.795 50.755 ;
        RECT 122.805 49.945 126.475 50.755 ;
        RECT 126.630 50.075 128.465 50.755 ;
        RECT 127.535 49.845 128.465 50.075 ;
        RECT 128.785 49.945 131.535 50.755 ;
        RECT 132.005 50.075 135.215 50.755 ;
        RECT 135.370 50.075 137.205 50.755 ;
        RECT 134.080 49.845 135.215 50.075 ;
        RECT 136.275 49.845 137.205 50.075 ;
        RECT 137.525 49.945 141.195 50.755 ;
        RECT 141.205 49.945 142.575 50.755 ;
        RECT 142.595 49.885 143.025 50.670 ;
        RECT 143.045 49.945 145.795 50.755 ;
        RECT 146.265 50.075 150.680 50.755 ;
        RECT 146.265 49.845 150.195 50.075 ;
        RECT 150.865 49.945 152.235 50.755 ;
      LAYER nwell ;
        RECT 90.870 46.725 152.430 49.555 ;
      LAYER pwell ;
        RECT 91.065 45.525 92.435 46.335 ;
        RECT 97.415 46.205 98.345 46.425 ;
        RECT 101.175 46.205 102.515 46.435 ;
        RECT 92.905 45.525 102.515 46.205 ;
        RECT 102.565 45.525 103.935 46.335 ;
        RECT 103.955 45.610 104.385 46.395 ;
        RECT 105.325 46.235 106.255 46.435 ;
        RECT 107.585 46.235 108.535 46.435 ;
        RECT 105.325 45.755 108.535 46.235 ;
        RECT 117.745 46.205 118.665 46.435 ;
        RECT 121.495 46.205 122.425 46.425 ;
        RECT 105.470 45.555 108.535 45.755 ;
        RECT 91.205 45.315 91.375 45.525 ;
        RECT 92.585 45.475 92.755 45.505 ;
        RECT 92.580 45.365 92.755 45.475 ;
        RECT 92.585 45.315 92.755 45.365 ;
        RECT 93.045 45.335 93.215 45.525 ;
        RECT 96.270 45.315 96.440 45.505 ;
        RECT 99.020 45.365 99.140 45.475 ;
        RECT 91.065 44.505 92.435 45.315 ;
        RECT 92.445 44.505 96.115 45.315 ;
        RECT 96.125 44.405 98.735 45.315 ;
        RECT 99.345 45.285 100.280 45.315 ;
        RECT 102.240 45.285 102.410 45.505 ;
        RECT 102.705 45.315 102.875 45.525 ;
        RECT 104.555 45.370 104.715 45.480 ;
        RECT 105.470 45.335 105.640 45.555 ;
        RECT 107.600 45.525 108.535 45.555 ;
        RECT 108.630 45.525 117.735 46.205 ;
        RECT 117.745 45.525 126.935 46.205 ;
        RECT 126.955 45.525 128.305 46.435 ;
        RECT 128.325 45.525 129.695 46.335 ;
        RECT 129.715 45.610 130.145 46.395 ;
        RECT 130.165 45.525 135.675 46.335 ;
        RECT 135.685 45.525 141.195 46.335 ;
        RECT 141.205 45.525 146.715 46.335 ;
        RECT 146.725 45.525 150.395 46.335 ;
        RECT 150.865 45.525 152.235 46.335 ;
        RECT 106.385 45.335 106.555 45.505 ;
        RECT 106.385 45.315 106.550 45.335 ;
        RECT 106.845 45.315 107.015 45.505 ;
        RECT 113.285 45.315 113.455 45.505 ;
        RECT 114.665 45.315 114.835 45.505 ;
        RECT 115.125 45.315 115.295 45.505 ;
        RECT 117.425 45.315 117.595 45.525 ;
        RECT 121.105 45.315 121.275 45.505 ;
        RECT 122.485 45.315 122.655 45.505 ;
        RECT 126.625 45.335 126.795 45.525 ;
        RECT 127.085 45.335 127.255 45.525 ;
        RECT 128.465 45.335 128.635 45.525 ;
        RECT 129.380 45.315 129.550 45.505 ;
        RECT 129.845 45.315 130.015 45.505 ;
        RECT 130.305 45.335 130.475 45.525 ;
        RECT 132.145 45.315 132.315 45.505 ;
        RECT 132.615 45.360 132.775 45.470 ;
        RECT 134.445 45.315 134.615 45.505 ;
        RECT 134.905 45.315 135.075 45.505 ;
        RECT 135.825 45.335 135.995 45.525 ;
        RECT 136.740 45.315 136.910 45.505 ;
        RECT 138.125 45.335 138.295 45.505 ;
        RECT 138.130 45.315 138.295 45.335 ;
        RECT 140.425 45.315 140.595 45.505 ;
        RECT 141.345 45.335 141.515 45.525 ;
        RECT 144.105 45.315 144.275 45.505 ;
        RECT 144.565 45.315 144.735 45.505 ;
        RECT 146.405 45.315 146.575 45.505 ;
        RECT 146.865 45.335 147.035 45.525 ;
        RECT 147.785 45.315 147.955 45.505 ;
        RECT 150.540 45.365 150.660 45.475 ;
        RECT 151.925 45.315 152.095 45.525 ;
        RECT 99.345 45.085 102.410 45.285 ;
        RECT 99.345 44.605 102.555 45.085 ;
        RECT 99.345 44.405 100.295 44.605 ;
        RECT 101.625 44.405 102.555 44.605 ;
        RECT 102.565 44.505 104.395 45.315 ;
        RECT 104.715 44.635 106.550 45.315 ;
        RECT 104.715 44.405 105.645 44.635 ;
        RECT 106.705 44.505 110.375 45.315 ;
        RECT 110.385 44.635 113.595 45.315 ;
        RECT 110.385 44.405 111.520 44.635 ;
        RECT 113.615 44.405 114.965 45.315 ;
        RECT 114.985 44.505 116.815 45.315 ;
        RECT 116.835 44.445 117.265 45.230 ;
        RECT 117.285 44.505 120.955 45.315 ;
        RECT 120.965 44.505 122.335 45.315 ;
        RECT 122.455 44.635 125.920 45.315 ;
        RECT 125.000 44.405 125.920 44.635 ;
        RECT 126.025 44.405 129.695 45.315 ;
        RECT 129.705 44.505 131.075 45.315 ;
        RECT 131.095 44.405 132.445 45.315 ;
        RECT 133.395 44.405 134.745 45.315 ;
        RECT 134.765 44.505 136.595 45.315 ;
        RECT 136.625 44.405 137.975 45.315 ;
        RECT 138.130 44.635 139.965 45.315 ;
        RECT 140.285 44.635 142.575 45.315 ;
        RECT 139.035 44.405 139.965 44.635 ;
        RECT 141.655 44.405 142.575 44.635 ;
        RECT 142.595 44.445 143.025 45.230 ;
        RECT 143.045 44.535 144.415 45.315 ;
        RECT 144.425 44.505 146.255 45.315 ;
        RECT 146.275 44.405 147.625 45.315 ;
        RECT 147.645 44.505 150.395 45.315 ;
        RECT 150.865 44.505 152.235 45.315 ;
      LAYER nwell ;
        RECT 90.870 41.285 152.430 44.115 ;
      LAYER pwell ;
        RECT 91.065 40.085 92.435 40.895 ;
        RECT 92.445 40.085 93.815 40.865 ;
        RECT 93.825 40.085 97.495 40.895 ;
        RECT 97.505 40.085 98.875 40.895 ;
        RECT 98.885 40.085 101.495 40.995 ;
        RECT 101.645 40.085 103.475 40.895 ;
        RECT 103.955 40.170 104.385 40.955 ;
        RECT 104.405 40.085 109.915 40.895 ;
        RECT 109.925 40.085 115.435 40.895 ;
        RECT 115.445 40.085 120.955 40.895 ;
        RECT 120.965 40.085 126.475 40.895 ;
        RECT 126.485 40.085 129.235 40.895 ;
        RECT 129.715 40.170 130.145 40.955 ;
        RECT 130.165 40.085 135.675 40.895 ;
        RECT 135.685 40.085 138.435 40.895 ;
        RECT 138.905 40.085 140.255 40.995 ;
        RECT 145.715 40.765 146.645 40.985 ;
        RECT 149.475 40.765 150.395 40.995 ;
        RECT 141.205 40.085 150.395 40.765 ;
        RECT 150.865 40.085 152.235 40.895 ;
        RECT 91.205 39.875 91.375 40.085 ;
        RECT 92.585 39.875 92.755 40.085 ;
        RECT 93.965 39.895 94.135 40.085 ;
        RECT 96.260 39.925 96.380 40.035 ;
        RECT 96.725 39.875 96.895 40.065 ;
        RECT 97.645 39.895 97.815 40.085 ;
        RECT 99.030 39.895 99.200 40.085 ;
        RECT 99.480 39.925 99.600 40.035 ;
        RECT 91.065 39.065 92.435 39.875 ;
        RECT 92.445 39.065 96.115 39.875 ;
        RECT 96.585 39.195 99.335 39.875 ;
        RECT 99.950 39.845 100.120 40.065 ;
        RECT 101.785 39.895 101.955 40.085 ;
        RECT 102.705 39.875 102.875 40.065 ;
        RECT 103.620 39.925 103.740 40.035 ;
        RECT 104.085 39.875 104.255 40.065 ;
        RECT 104.545 39.895 104.715 40.085 ;
        RECT 106.845 39.875 107.015 40.065 ;
        RECT 110.065 39.895 110.235 40.085 ;
        RECT 110.985 39.875 111.155 40.065 ;
        RECT 113.745 39.875 113.915 40.065 ;
        RECT 114.210 39.875 114.380 40.065 ;
        RECT 115.585 39.895 115.755 40.085 ;
        RECT 116.055 39.920 116.215 40.030 ;
        RECT 117.425 39.875 117.595 40.065 ;
        RECT 119.265 39.875 119.435 40.065 ;
        RECT 121.105 39.895 121.275 40.085 ;
        RECT 122.485 39.875 122.655 40.065 ;
        RECT 125.705 39.875 125.875 40.065 ;
        RECT 126.625 39.895 126.795 40.085 ;
        RECT 129.380 39.925 129.500 40.035 ;
        RECT 130.305 39.895 130.475 40.085 ;
        RECT 131.225 39.875 131.395 40.065 ;
        RECT 132.605 39.875 132.775 40.065 ;
        RECT 133.065 39.875 133.235 40.065 ;
        RECT 135.825 40.035 135.995 40.085 ;
        RECT 135.820 39.925 135.995 40.035 ;
        RECT 135.825 39.895 135.995 39.925 ;
        RECT 136.290 39.875 136.460 40.065 ;
        RECT 138.580 39.925 138.700 40.035 ;
        RECT 139.050 39.895 139.220 40.085 ;
        RECT 140.435 39.930 140.595 40.040 ;
        RECT 141.345 39.875 141.515 40.085 ;
        RECT 141.815 39.920 141.975 40.030 ;
        RECT 143.185 39.875 143.355 40.065 ;
        RECT 150.545 40.035 150.715 40.065 ;
        RECT 146.415 39.920 146.575 40.030 ;
        RECT 150.540 39.925 150.715 40.035 ;
        RECT 150.545 39.875 150.715 39.925 ;
        RECT 151.925 39.875 152.095 40.085 ;
        RECT 101.610 39.845 102.555 39.875 ;
        RECT 98.405 38.965 99.335 39.195 ;
        RECT 99.805 39.165 102.555 39.845 ;
        RECT 101.610 38.965 102.555 39.165 ;
        RECT 102.565 39.065 103.935 39.875 ;
        RECT 103.945 39.195 106.695 39.875 ;
        RECT 105.765 38.965 106.695 39.195 ;
        RECT 106.705 39.065 108.075 39.875 ;
        RECT 108.085 38.965 111.295 39.875 ;
        RECT 111.305 39.195 114.055 39.875 ;
        RECT 111.305 38.965 112.235 39.195 ;
        RECT 114.065 38.965 115.895 39.875 ;
        RECT 116.835 39.005 117.265 39.790 ;
        RECT 117.285 39.065 119.115 39.875 ;
        RECT 119.205 38.965 122.205 39.875 ;
        RECT 122.345 38.965 125.555 39.875 ;
        RECT 125.565 38.965 128.775 39.875 ;
        RECT 128.785 39.645 131.395 39.875 ;
        RECT 128.785 38.965 131.535 39.645 ;
        RECT 131.555 38.965 132.905 39.875 ;
        RECT 132.925 39.065 135.675 39.875 ;
        RECT 136.145 38.965 139.795 39.875 ;
        RECT 139.825 38.965 141.640 39.875 ;
        RECT 142.595 39.005 143.025 39.790 ;
        RECT 143.085 38.965 146.255 39.875 ;
        RECT 147.280 39.195 150.745 39.875 ;
        RECT 147.280 38.965 148.200 39.195 ;
        RECT 150.865 39.065 152.235 39.875 ;
      LAYER nwell ;
        RECT 90.870 35.845 152.430 38.675 ;
      LAYER pwell ;
        RECT 91.065 34.645 92.435 35.455 ;
        RECT 94.250 35.355 95.195 35.555 ;
        RECT 92.445 34.675 95.195 35.355 ;
        RECT 95.205 35.355 96.135 35.555 ;
        RECT 97.465 35.355 98.415 35.555 ;
        RECT 95.205 34.875 98.415 35.355 ;
        RECT 91.205 34.435 91.375 34.645 ;
        RECT 92.590 34.625 92.760 34.675 ;
        RECT 94.250 34.645 95.195 34.675 ;
        RECT 95.350 34.675 98.415 34.875 ;
        RECT 92.585 34.455 92.760 34.625 ;
        RECT 95.350 34.455 95.520 34.675 ;
        RECT 97.480 34.645 98.415 34.675 ;
        RECT 98.425 34.645 102.555 35.555 ;
        RECT 102.575 34.645 103.925 35.555 ;
        RECT 103.955 34.730 104.385 35.515 ;
        RECT 104.555 34.645 108.210 35.555 ;
        RECT 109.615 34.645 113.270 35.555 ;
        RECT 113.615 34.645 114.965 35.555 ;
        RECT 114.985 34.645 118.195 35.555 ;
        RECT 118.205 34.645 120.035 35.455 ;
        RECT 121.850 35.355 122.795 35.555 ;
        RECT 120.045 34.675 122.795 35.355 ;
        RECT 92.585 34.435 92.755 34.455 ;
        RECT 91.065 33.625 92.435 34.435 ;
        RECT 92.445 33.625 97.955 34.435 ;
        RECT 98.110 34.405 98.280 34.625 ;
        RECT 102.245 34.455 102.415 34.645 ;
        RECT 102.705 34.455 102.875 34.645 ;
        RECT 104.555 34.625 104.715 34.645 ;
        RECT 109.615 34.625 109.775 34.645 ;
        RECT 99.770 34.405 100.715 34.435 ;
        RECT 97.965 33.725 100.715 34.405 ;
        RECT 99.770 33.525 100.715 33.725 ;
        RECT 100.725 34.405 101.670 34.435 ;
        RECT 103.160 34.405 103.330 34.625 ;
        RECT 103.620 34.485 103.740 34.595 ;
        RECT 104.085 34.435 104.255 34.625 ;
        RECT 104.545 34.455 104.715 34.625 ;
        RECT 108.695 34.490 108.855 34.600 ;
        RECT 109.605 34.455 109.775 34.625 ;
        RECT 110.065 34.435 110.235 34.625 ;
        RECT 110.520 34.485 110.640 34.595 ;
        RECT 110.985 34.435 111.155 34.625 ;
        RECT 114.665 34.455 114.835 34.645 ;
        RECT 115.125 34.455 115.295 34.645 ;
        RECT 116.045 34.455 116.215 34.625 ;
        RECT 116.500 34.485 116.620 34.595 ;
        RECT 117.420 34.485 117.540 34.595 ;
        RECT 116.045 34.435 116.210 34.455 ;
        RECT 100.725 33.725 103.475 34.405 ;
        RECT 100.725 33.525 101.670 33.725 ;
        RECT 103.945 33.525 107.615 34.435 ;
        RECT 107.625 33.755 110.375 34.435 ;
        RECT 107.625 33.525 108.555 33.755 ;
        RECT 110.845 33.525 114.055 34.435 ;
        RECT 114.375 33.755 116.210 34.435 ;
        RECT 117.890 34.405 118.060 34.625 ;
        RECT 118.345 34.455 118.515 34.645 ;
        RECT 120.190 34.455 120.360 34.675 ;
        RECT 121.850 34.645 122.795 34.675 ;
        RECT 122.805 35.325 123.730 35.555 ;
        RECT 122.805 34.645 126.475 35.325 ;
        RECT 126.485 34.645 129.695 35.555 ;
        RECT 129.715 34.730 130.145 35.515 ;
        RECT 130.165 34.645 133.375 35.555 ;
        RECT 133.385 34.645 137.040 35.555 ;
        RECT 137.545 34.645 138.895 35.555 ;
        RECT 139.835 34.645 141.185 35.555 ;
        RECT 145.715 35.325 146.645 35.545 ;
        RECT 149.475 35.325 150.395 35.555 ;
        RECT 141.205 34.645 150.395 35.325 ;
        RECT 150.865 34.645 152.235 35.455 ;
        RECT 120.655 34.480 120.815 34.590 ;
        RECT 122.485 34.435 122.655 34.625 ;
        RECT 122.950 34.455 123.120 34.645 ;
        RECT 125.245 34.435 125.415 34.625 ;
        RECT 125.715 34.480 125.875 34.590 ;
        RECT 126.625 34.435 126.795 34.625 ;
        RECT 129.385 34.455 129.555 34.645 ;
        RECT 129.845 34.435 130.015 34.625 ;
        RECT 130.305 34.455 130.475 34.645 ;
        RECT 133.530 34.455 133.700 34.645 ;
        RECT 133.985 34.435 134.155 34.625 ;
        RECT 134.445 34.435 134.615 34.625 ;
        RECT 137.200 34.485 137.320 34.595 ;
        RECT 138.580 34.455 138.750 34.645 ;
        RECT 139.055 34.490 139.215 34.600 ;
        RECT 139.965 34.435 140.135 34.645 ;
        RECT 141.345 34.455 141.515 34.645 ;
        RECT 143.185 34.435 143.355 34.625 ;
        RECT 145.940 34.485 146.060 34.595 ;
        RECT 146.410 34.435 146.580 34.625 ;
        RECT 147.785 34.435 147.955 34.625 ;
        RECT 149.160 34.485 149.280 34.595 ;
        RECT 150.535 34.435 150.705 34.625 ;
        RECT 151.925 34.435 152.095 34.645 ;
        RECT 119.550 34.405 120.495 34.435 ;
        RECT 114.375 33.525 115.305 33.755 ;
        RECT 116.835 33.565 117.265 34.350 ;
        RECT 117.745 33.725 120.495 34.405 ;
        RECT 119.550 33.525 120.495 33.725 ;
        RECT 121.435 33.525 122.785 34.435 ;
        RECT 122.815 33.525 125.545 34.435 ;
        RECT 126.485 33.525 129.695 34.435 ;
        RECT 129.705 33.625 131.075 34.435 ;
        RECT 131.085 33.525 134.295 34.435 ;
        RECT 134.305 33.625 139.815 34.435 ;
        RECT 139.825 33.625 142.575 34.435 ;
        RECT 142.595 33.565 143.025 34.350 ;
        RECT 143.045 33.625 145.795 34.435 ;
        RECT 146.265 33.525 147.615 34.435 ;
        RECT 147.655 33.525 149.005 34.435 ;
        RECT 149.485 33.655 150.855 34.435 ;
        RECT 150.865 33.625 152.235 34.435 ;
      LAYER nwell ;
        RECT 90.870 30.405 152.430 33.235 ;
      LAYER pwell ;
        RECT 91.065 29.205 92.435 30.015 ;
        RECT 92.445 29.205 93.815 29.985 ;
        RECT 93.825 29.205 97.495 30.015 ;
        RECT 98.425 29.205 99.795 29.985 ;
        RECT 99.805 29.205 103.475 30.015 ;
        RECT 103.955 29.290 104.385 30.075 ;
        RECT 104.405 29.205 106.235 30.015 ;
        RECT 106.245 29.205 107.615 29.985 ;
        RECT 107.625 29.205 113.135 30.015 ;
        RECT 114.065 29.205 115.435 29.985 ;
        RECT 115.445 29.205 116.815 30.015 ;
        RECT 116.835 29.290 117.265 30.075 ;
        RECT 117.285 29.205 118.655 30.015 ;
        RECT 118.675 29.205 120.025 30.115 ;
        RECT 120.045 29.205 121.875 30.015 ;
        RECT 121.885 29.205 123.255 29.985 ;
        RECT 123.265 29.205 128.775 30.015 ;
        RECT 129.715 29.290 130.145 30.075 ;
        RECT 130.165 29.205 131.535 29.985 ;
        RECT 131.545 29.205 137.055 30.015 ;
        RECT 137.525 29.205 138.895 29.985 ;
        RECT 138.905 29.205 142.575 30.015 ;
        RECT 142.595 29.290 143.025 30.075 ;
        RECT 143.705 29.885 147.635 30.115 ;
        RECT 143.220 29.205 147.635 29.885 ;
        RECT 147.645 29.205 149.015 30.015 ;
        RECT 149.025 29.205 150.855 29.885 ;
        RECT 150.865 29.205 152.235 30.015 ;
        RECT 91.205 29.015 91.375 29.205 ;
        RECT 92.595 29.015 92.765 29.205 ;
        RECT 93.965 29.015 94.135 29.205 ;
        RECT 97.655 29.050 97.815 29.160 ;
        RECT 98.575 29.015 98.745 29.205 ;
        RECT 99.945 29.015 100.115 29.205 ;
        RECT 103.620 29.045 103.740 29.155 ;
        RECT 104.545 29.015 104.715 29.205 ;
        RECT 106.395 29.015 106.565 29.205 ;
        RECT 107.765 29.015 107.935 29.205 ;
        RECT 113.295 29.050 113.455 29.160 ;
        RECT 114.215 29.015 114.385 29.205 ;
        RECT 115.585 29.015 115.755 29.205 ;
        RECT 117.425 29.015 117.595 29.205 ;
        RECT 119.725 29.015 119.895 29.205 ;
        RECT 120.185 29.015 120.355 29.205 ;
        RECT 122.935 29.015 123.105 29.205 ;
        RECT 123.405 29.015 123.575 29.205 ;
        RECT 128.935 29.050 129.095 29.160 ;
        RECT 131.215 29.015 131.385 29.205 ;
        RECT 131.685 29.015 131.855 29.205 ;
        RECT 137.200 29.045 137.320 29.155 ;
        RECT 138.575 29.015 138.745 29.205 ;
        RECT 139.045 29.015 139.215 29.205 ;
        RECT 143.220 29.185 143.330 29.205 ;
        RECT 143.160 29.015 143.330 29.185 ;
        RECT 147.785 29.015 147.955 29.205 ;
        RECT 150.545 29.015 150.715 29.205 ;
        RECT 151.925 29.015 152.095 29.205 ;
      LAYER li1 ;
        RECT 71.250 194.345 119.550 194.515 ;
        RECT 71.335 193.255 72.545 194.345 ;
        RECT 72.715 193.910 78.060 194.345 ;
        RECT 71.335 192.545 71.855 193.085 ;
        RECT 72.025 192.715 72.545 193.255 ;
        RECT 71.335 191.795 72.545 192.545 ;
        RECT 74.300 192.340 74.640 193.170 ;
        RECT 76.120 192.660 76.470 193.910 ;
        RECT 78.235 193.255 80.825 194.345 ;
        RECT 78.235 192.565 79.445 193.085 ;
        RECT 79.615 192.735 80.825 193.255 ;
        RECT 80.995 193.375 81.305 194.175 ;
        RECT 81.475 193.545 81.785 194.345 ;
        RECT 81.955 193.715 82.215 194.175 ;
        RECT 82.385 193.885 82.640 194.345 ;
        RECT 82.815 193.715 83.075 194.175 ;
        RECT 81.955 193.545 83.075 193.715 ;
        RECT 80.995 193.205 82.025 193.375 ;
        RECT 72.715 191.795 78.060 192.340 ;
        RECT 78.235 191.795 80.825 192.565 ;
        RECT 80.995 192.295 81.165 193.205 ;
        RECT 81.335 192.465 81.685 193.035 ;
        RECT 81.855 192.955 82.025 193.205 ;
        RECT 82.815 193.295 83.075 193.545 ;
        RECT 83.245 193.475 83.530 194.345 ;
        RECT 82.815 193.125 83.570 193.295 ;
        RECT 84.215 193.180 84.505 194.345 ;
        RECT 84.675 193.255 85.885 194.345 ;
        RECT 81.855 192.785 82.995 192.955 ;
        RECT 83.165 192.615 83.570 193.125 ;
        RECT 81.920 192.445 83.570 192.615 ;
        RECT 84.675 192.545 85.195 193.085 ;
        RECT 85.365 192.715 85.885 193.255 ;
        RECT 86.055 193.205 86.440 194.175 ;
        RECT 86.610 193.885 86.935 194.345 ;
        RECT 87.455 193.715 87.735 194.175 ;
        RECT 86.610 193.495 87.735 193.715 ;
        RECT 80.995 191.965 81.295 192.295 ;
        RECT 81.465 191.795 81.740 192.275 ;
        RECT 81.920 192.055 82.215 192.445 ;
        RECT 82.385 191.795 82.640 192.275 ;
        RECT 82.815 192.055 83.075 192.445 ;
        RECT 83.245 191.795 83.525 192.275 ;
        RECT 84.215 191.795 84.505 192.520 ;
        RECT 84.675 191.795 85.885 192.545 ;
        RECT 86.055 192.535 86.335 193.205 ;
        RECT 86.610 193.035 87.060 193.495 ;
        RECT 87.925 193.325 88.325 194.175 ;
        RECT 88.725 193.885 88.995 194.345 ;
        RECT 89.165 193.715 89.450 194.175 ;
        RECT 89.735 193.910 95.080 194.345 ;
        RECT 86.505 192.705 87.060 193.035 ;
        RECT 87.230 192.765 88.325 193.325 ;
        RECT 86.610 192.595 87.060 192.705 ;
        RECT 86.055 191.965 86.440 192.535 ;
        RECT 86.610 192.425 87.735 192.595 ;
        RECT 86.610 191.795 86.935 192.255 ;
        RECT 87.455 191.965 87.735 192.425 ;
        RECT 87.925 191.965 88.325 192.765 ;
        RECT 88.495 193.495 89.450 193.715 ;
        RECT 88.495 192.595 88.705 193.495 ;
        RECT 88.875 192.765 89.565 193.325 ;
        RECT 88.495 192.425 89.450 192.595 ;
        RECT 88.725 191.795 88.995 192.255 ;
        RECT 89.165 191.965 89.450 192.425 ;
        RECT 91.320 192.340 91.660 193.170 ;
        RECT 93.140 192.660 93.490 193.910 ;
        RECT 95.255 193.255 96.925 194.345 ;
        RECT 95.255 192.565 96.005 193.085 ;
        RECT 96.175 192.735 96.925 193.255 ;
        RECT 97.095 193.180 97.385 194.345 ;
        RECT 97.555 193.255 100.145 194.345 ;
        RECT 97.555 192.565 98.765 193.085 ;
        RECT 98.935 192.735 100.145 193.255 ;
        RECT 100.500 193.375 100.890 193.550 ;
        RECT 101.375 193.545 101.705 194.345 ;
        RECT 101.875 193.555 102.410 194.175 ;
        RECT 102.615 193.910 107.960 194.345 ;
        RECT 100.500 193.205 101.925 193.375 ;
        RECT 89.735 191.795 95.080 192.340 ;
        RECT 95.255 191.795 96.925 192.565 ;
        RECT 97.095 191.795 97.385 192.520 ;
        RECT 97.555 191.795 100.145 192.565 ;
        RECT 100.375 192.475 100.730 193.035 ;
        RECT 100.900 192.305 101.070 193.205 ;
        RECT 101.240 192.475 101.505 193.035 ;
        RECT 101.755 192.705 101.925 193.205 ;
        RECT 102.095 192.535 102.410 193.555 ;
        RECT 100.480 191.795 100.720 192.305 ;
        RECT 100.900 191.975 101.180 192.305 ;
        RECT 101.410 191.795 101.625 192.305 ;
        RECT 101.795 191.965 102.410 192.535 ;
        RECT 104.200 192.340 104.540 193.170 ;
        RECT 106.020 192.660 106.370 193.910 ;
        RECT 108.135 193.255 109.805 194.345 ;
        RECT 108.135 192.565 108.885 193.085 ;
        RECT 109.055 192.735 109.805 193.255 ;
        RECT 109.975 193.180 110.265 194.345 ;
        RECT 110.895 193.375 111.205 194.175 ;
        RECT 111.375 193.545 111.685 194.345 ;
        RECT 111.855 193.715 112.115 194.175 ;
        RECT 112.285 193.885 112.540 194.345 ;
        RECT 112.715 193.715 112.975 194.175 ;
        RECT 111.855 193.545 112.975 193.715 ;
        RECT 110.895 193.205 111.925 193.375 ;
        RECT 102.615 191.795 107.960 192.340 ;
        RECT 108.135 191.795 109.805 192.565 ;
        RECT 109.975 191.795 110.265 192.520 ;
        RECT 110.895 192.295 111.065 193.205 ;
        RECT 111.235 192.465 111.585 193.035 ;
        RECT 111.755 192.955 111.925 193.205 ;
        RECT 112.715 193.295 112.975 193.545 ;
        RECT 113.145 193.475 113.430 194.345 ;
        RECT 112.715 193.125 113.470 193.295 ;
        RECT 113.655 193.255 117.165 194.345 ;
        RECT 111.755 192.785 112.895 192.955 ;
        RECT 113.065 192.615 113.470 193.125 ;
        RECT 111.820 192.445 113.470 192.615 ;
        RECT 113.655 192.565 115.305 193.085 ;
        RECT 115.475 192.735 117.165 193.255 ;
        RECT 118.255 193.255 119.465 194.345 ;
        RECT 118.255 192.715 118.775 193.255 ;
        RECT 110.895 191.965 111.195 192.295 ;
        RECT 111.365 191.795 111.640 192.275 ;
        RECT 111.820 192.055 112.115 192.445 ;
        RECT 112.285 191.795 112.540 192.275 ;
        RECT 112.715 192.055 112.975 192.445 ;
        RECT 113.145 191.795 113.425 192.275 ;
        RECT 113.655 191.795 117.165 192.565 ;
        RECT 118.945 192.545 119.465 193.085 ;
        RECT 118.255 191.795 119.465 192.545 ;
        RECT 71.250 191.625 119.550 191.795 ;
        RECT 71.335 190.875 72.545 191.625 ;
        RECT 72.805 191.075 72.975 191.455 ;
        RECT 73.155 191.245 73.485 191.625 ;
        RECT 72.805 190.905 73.470 191.075 ;
        RECT 73.665 190.950 73.925 191.455 ;
        RECT 71.335 190.335 71.855 190.875 ;
        RECT 72.025 190.165 72.545 190.705 ;
        RECT 72.735 190.355 73.065 190.725 ;
        RECT 73.300 190.650 73.470 190.905 ;
        RECT 73.300 190.320 73.585 190.650 ;
        RECT 73.300 190.175 73.470 190.320 ;
        RECT 71.335 189.075 72.545 190.165 ;
        RECT 72.805 190.005 73.470 190.175 ;
        RECT 73.755 190.150 73.925 190.950 ;
        RECT 74.095 190.855 76.685 191.625 ;
        RECT 77.315 190.965 77.575 191.295 ;
        RECT 77.770 190.995 77.995 191.625 ;
        RECT 78.210 190.990 78.455 191.450 ;
        RECT 78.705 191.165 78.975 191.625 ;
        RECT 79.145 191.175 79.985 191.345 ;
        RECT 80.545 191.265 80.875 191.625 ;
        RECT 74.095 190.335 75.305 190.855 ;
        RECT 75.475 190.165 76.685 190.685 ;
        RECT 72.805 189.245 72.975 190.005 ;
        RECT 73.155 189.075 73.485 189.835 ;
        RECT 73.655 189.245 73.925 190.150 ;
        RECT 74.095 189.075 76.685 190.165 ;
        RECT 77.315 190.040 77.485 190.965 ;
        RECT 78.210 190.715 78.380 190.990 ;
        RECT 79.145 190.715 79.315 191.175 ;
        RECT 81.045 191.095 81.240 191.365 ;
        RECT 77.655 190.385 78.380 190.715 ;
        RECT 78.550 190.385 79.315 190.715 ;
        RECT 78.210 190.175 78.380 190.385 ;
        RECT 79.105 190.260 79.315 190.385 ;
        RECT 79.485 190.670 80.190 190.975 ;
        RECT 80.635 190.945 81.240 191.095 ;
        RECT 80.430 190.925 81.240 190.945 ;
        RECT 77.315 189.255 77.575 190.040 ;
        RECT 77.745 189.075 78.030 190.140 ;
        RECT 78.210 189.845 78.935 190.175 ;
        RECT 78.210 189.275 78.455 189.845 ;
        RECT 79.105 189.700 79.295 190.260 ;
        RECT 79.485 190.150 79.800 190.670 ;
        RECT 80.430 190.475 80.805 190.925 ;
        RECT 79.465 189.800 79.800 190.150 ;
        RECT 79.970 189.705 80.305 190.355 ;
        RECT 80.635 190.215 80.805 190.475 ;
        RECT 80.985 190.385 81.315 190.755 ;
        RECT 80.635 190.045 81.320 190.215 ;
        RECT 79.105 189.675 79.320 189.700 ;
        RECT 79.105 189.665 79.345 189.675 ;
        RECT 79.105 189.645 79.360 189.665 ;
        RECT 79.120 189.625 79.360 189.645 ;
        RECT 79.130 189.620 79.360 189.625 ;
        RECT 79.130 189.605 79.455 189.620 ;
        RECT 78.655 189.075 78.975 189.535 ;
        RECT 79.145 189.455 79.455 189.605 ;
        RECT 79.145 189.285 80.005 189.455 ;
        RECT 80.505 189.075 80.795 189.875 ;
        RECT 80.965 189.295 81.320 190.045 ;
        RECT 81.565 190.025 81.735 191.365 ;
        RECT 81.905 191.245 82.235 191.625 ;
        RECT 82.405 191.075 82.575 191.365 ;
        RECT 81.970 190.905 82.575 191.075 ;
        RECT 81.970 190.640 82.140 190.905 ;
        RECT 82.835 190.825 83.145 191.625 ;
        RECT 83.350 190.825 84.045 191.455 ;
        RECT 84.215 190.855 86.805 191.625 ;
        RECT 87.025 190.970 87.355 191.405 ;
        RECT 87.525 191.015 87.695 191.625 ;
        RECT 86.975 190.885 87.355 190.970 ;
        RECT 87.865 190.885 88.195 191.410 ;
        RECT 88.455 191.095 88.665 191.625 ;
        RECT 88.940 191.175 89.725 191.345 ;
        RECT 89.895 191.175 90.300 191.345 ;
        RECT 81.910 190.310 82.140 190.640 ;
        RECT 81.510 189.245 81.735 190.025 ;
        RECT 81.970 189.915 82.140 190.310 ;
        RECT 82.420 190.085 82.665 190.725 ;
        RECT 82.845 190.385 83.180 190.655 ;
        RECT 83.350 190.225 83.520 190.825 ;
        RECT 83.690 190.385 84.025 190.635 ;
        RECT 84.215 190.335 85.425 190.855 ;
        RECT 86.975 190.845 87.200 190.885 ;
        RECT 81.970 189.745 82.575 189.915 ;
        RECT 81.905 189.075 82.235 189.575 ;
        RECT 82.405 189.245 82.575 189.745 ;
        RECT 82.835 189.075 83.115 190.215 ;
        RECT 83.285 189.245 83.615 190.225 ;
        RECT 83.785 189.075 84.045 190.215 ;
        RECT 85.595 190.165 86.805 190.685 ;
        RECT 84.215 189.075 86.805 190.165 ;
        RECT 86.975 190.265 87.145 190.845 ;
        RECT 87.865 190.715 88.065 190.885 ;
        RECT 88.940 190.715 89.110 191.175 ;
        RECT 87.315 190.385 88.065 190.715 ;
        RECT 88.235 190.385 89.110 190.715 ;
        RECT 86.975 190.215 87.190 190.265 ;
        RECT 86.975 190.135 87.365 190.215 ;
        RECT 87.035 189.290 87.365 190.135 ;
        RECT 87.875 190.180 88.065 190.385 ;
        RECT 87.535 189.075 87.705 190.085 ;
        RECT 87.875 189.805 88.770 190.180 ;
        RECT 87.875 189.245 88.215 189.805 ;
        RECT 88.445 189.075 88.760 189.575 ;
        RECT 88.940 189.545 89.110 190.385 ;
        RECT 89.280 190.675 89.745 191.005 ;
        RECT 90.130 190.945 90.300 191.175 ;
        RECT 90.480 191.125 90.850 191.625 ;
        RECT 91.170 191.175 91.845 191.345 ;
        RECT 92.040 191.175 92.375 191.345 ;
        RECT 89.280 189.715 89.600 190.675 ;
        RECT 90.130 190.645 90.960 190.945 ;
        RECT 89.770 189.745 89.960 190.465 ;
        RECT 90.130 189.575 90.300 190.645 ;
        RECT 90.760 190.615 90.960 190.645 ;
        RECT 90.470 190.395 90.640 190.465 ;
        RECT 91.170 190.395 91.340 191.175 ;
        RECT 92.205 191.035 92.375 191.175 ;
        RECT 92.545 191.165 92.795 191.625 ;
        RECT 90.470 190.225 91.340 190.395 ;
        RECT 91.510 190.755 92.035 190.975 ;
        RECT 92.205 190.905 92.430 191.035 ;
        RECT 90.470 190.135 90.980 190.225 ;
        RECT 88.940 189.375 89.825 189.545 ;
        RECT 90.050 189.245 90.300 189.575 ;
        RECT 90.470 189.075 90.640 189.875 ;
        RECT 90.810 189.520 90.980 190.135 ;
        RECT 91.510 190.055 91.680 190.755 ;
        RECT 91.150 189.690 91.680 190.055 ;
        RECT 91.850 189.990 92.090 190.585 ;
        RECT 92.260 189.800 92.430 190.905 ;
        RECT 92.600 190.045 92.880 190.995 ;
        RECT 92.125 189.670 92.430 189.800 ;
        RECT 90.810 189.350 91.915 189.520 ;
        RECT 92.125 189.245 92.375 189.670 ;
        RECT 92.545 189.075 92.810 189.535 ;
        RECT 93.050 189.245 93.235 191.365 ;
        RECT 93.405 191.245 93.735 191.625 ;
        RECT 93.905 191.075 94.075 191.365 ;
        RECT 93.410 190.905 94.075 191.075 ;
        RECT 94.425 190.945 94.595 191.320 ;
        RECT 93.410 189.915 93.640 190.905 ;
        RECT 94.395 190.775 94.595 190.945 ;
        RECT 94.785 191.095 95.015 191.400 ;
        RECT 95.185 191.265 95.515 191.625 ;
        RECT 95.710 191.095 96.000 191.445 ;
        RECT 94.785 190.925 96.000 191.095 ;
        RECT 97.095 190.900 97.385 191.625 ;
        RECT 94.425 190.755 94.595 190.775 ;
        RECT 97.555 190.885 97.940 191.455 ;
        RECT 98.110 191.165 98.435 191.625 ;
        RECT 98.955 190.995 99.235 191.455 ;
        RECT 93.810 190.085 94.160 190.735 ;
        RECT 94.425 190.585 94.945 190.755 ;
        RECT 94.340 190.055 94.585 190.415 ;
        RECT 94.775 190.205 94.945 190.585 ;
        RECT 95.115 190.385 95.500 190.715 ;
        RECT 95.680 190.605 95.940 190.715 ;
        RECT 95.680 190.435 95.945 190.605 ;
        RECT 95.680 190.385 95.940 190.435 ;
        RECT 94.775 189.925 95.125 190.205 ;
        RECT 93.410 189.745 94.075 189.915 ;
        RECT 93.405 189.075 93.735 189.575 ;
        RECT 93.905 189.245 94.075 189.745 ;
        RECT 94.340 189.075 94.595 189.875 ;
        RECT 94.795 189.245 95.125 189.925 ;
        RECT 95.305 189.335 95.500 190.385 ;
        RECT 95.680 189.075 96.000 190.215 ;
        RECT 97.095 189.075 97.385 190.240 ;
        RECT 97.555 190.215 97.835 190.885 ;
        RECT 98.110 190.825 99.235 190.995 ;
        RECT 98.110 190.715 98.560 190.825 ;
        RECT 98.005 190.385 98.560 190.715 ;
        RECT 99.425 190.655 99.825 191.455 ;
        RECT 100.225 191.165 100.495 191.625 ;
        RECT 100.665 190.995 100.950 191.455 ;
        RECT 97.555 189.245 97.940 190.215 ;
        RECT 98.110 189.925 98.560 190.385 ;
        RECT 98.730 190.095 99.825 190.655 ;
        RECT 98.110 189.705 99.235 189.925 ;
        RECT 98.110 189.075 98.435 189.535 ;
        RECT 98.955 189.245 99.235 189.705 ;
        RECT 99.425 189.245 99.825 190.095 ;
        RECT 99.995 190.825 100.950 190.995 ;
        RECT 99.995 189.925 100.205 190.825 ;
        RECT 100.375 190.095 101.065 190.655 ;
        RECT 99.995 189.705 100.950 189.925 ;
        RECT 100.225 189.075 100.495 189.535 ;
        RECT 100.665 189.245 100.950 189.705 ;
        RECT 101.245 189.255 101.505 191.445 ;
        RECT 101.765 191.255 102.435 191.625 ;
        RECT 102.615 191.075 102.925 191.445 ;
        RECT 101.695 190.875 102.925 191.075 ;
        RECT 101.695 190.205 101.985 190.875 ;
        RECT 103.105 190.695 103.335 191.335 ;
        RECT 103.515 190.895 103.805 191.625 ;
        RECT 103.995 190.855 105.665 191.625 ;
        RECT 105.925 191.075 106.095 191.365 ;
        RECT 106.265 191.245 106.595 191.625 ;
        RECT 105.925 190.905 106.530 191.075 ;
        RECT 102.165 190.385 102.630 190.695 ;
        RECT 102.810 190.385 103.335 190.695 ;
        RECT 103.515 190.385 103.815 190.715 ;
        RECT 103.995 190.335 104.745 190.855 ;
        RECT 101.695 189.985 102.465 190.205 ;
        RECT 101.675 189.075 102.015 189.805 ;
        RECT 102.195 189.255 102.465 189.985 ;
        RECT 102.645 189.965 103.805 190.205 ;
        RECT 104.915 190.165 105.665 190.685 ;
        RECT 102.645 189.255 102.875 189.965 ;
        RECT 103.045 189.075 103.375 189.785 ;
        RECT 103.545 189.255 103.805 189.965 ;
        RECT 103.995 189.075 105.665 190.165 ;
        RECT 105.835 190.085 106.080 190.725 ;
        RECT 106.360 190.640 106.530 190.905 ;
        RECT 106.360 190.310 106.590 190.640 ;
        RECT 106.360 189.915 106.530 190.310 ;
        RECT 105.925 189.745 106.530 189.915 ;
        RECT 106.765 190.025 106.935 191.365 ;
        RECT 107.260 191.095 107.455 191.365 ;
        RECT 107.625 191.265 107.955 191.625 ;
        RECT 108.515 191.175 109.355 191.345 ;
        RECT 107.260 190.945 107.865 191.095 ;
        RECT 107.260 190.925 108.070 190.945 ;
        RECT 107.185 190.385 107.515 190.755 ;
        RECT 107.695 190.475 108.070 190.925 ;
        RECT 108.310 190.670 109.015 190.975 ;
        RECT 107.695 190.215 107.865 190.475 ;
        RECT 107.180 190.045 107.865 190.215 ;
        RECT 105.925 189.245 106.095 189.745 ;
        RECT 106.265 189.075 106.595 189.575 ;
        RECT 106.765 189.245 106.990 190.025 ;
        RECT 107.180 189.295 107.535 190.045 ;
        RECT 107.705 189.075 107.995 189.875 ;
        RECT 108.195 189.705 108.530 190.355 ;
        RECT 108.700 190.150 109.015 190.670 ;
        RECT 109.185 190.715 109.355 191.175 ;
        RECT 109.525 191.165 109.795 191.625 ;
        RECT 110.045 190.990 110.290 191.450 ;
        RECT 110.505 190.995 110.730 191.625 ;
        RECT 110.120 190.715 110.290 190.990 ;
        RECT 110.925 190.965 111.185 191.295 ;
        RECT 111.355 191.080 116.700 191.625 ;
        RECT 109.185 190.385 109.950 190.715 ;
        RECT 110.120 190.385 110.845 190.715 ;
        RECT 109.185 190.260 109.395 190.385 ;
        RECT 108.700 189.800 109.035 190.150 ;
        RECT 109.205 189.700 109.395 190.260 ;
        RECT 110.120 190.175 110.290 190.385 ;
        RECT 109.565 189.845 110.290 190.175 ;
        RECT 109.180 189.675 109.395 189.700 ;
        RECT 109.155 189.665 109.395 189.675 ;
        RECT 109.140 189.645 109.395 189.665 ;
        RECT 109.140 189.625 109.380 189.645 ;
        RECT 109.140 189.620 109.370 189.625 ;
        RECT 109.045 189.605 109.370 189.620 ;
        RECT 109.045 189.455 109.355 189.605 ;
        RECT 108.495 189.285 109.355 189.455 ;
        RECT 109.525 189.075 109.845 189.535 ;
        RECT 110.045 189.275 110.290 189.845 ;
        RECT 110.470 189.075 110.755 190.140 ;
        RECT 111.015 190.040 111.185 190.965 ;
        RECT 112.940 190.250 113.280 191.080 ;
        RECT 116.875 190.950 117.135 191.455 ;
        RECT 117.315 191.245 117.645 191.625 ;
        RECT 117.825 191.075 117.995 191.455 ;
        RECT 110.925 189.255 111.185 190.040 ;
        RECT 114.760 189.510 115.110 190.760 ;
        RECT 116.875 190.150 117.055 190.950 ;
        RECT 117.330 190.905 117.995 191.075 ;
        RECT 117.330 190.650 117.500 190.905 ;
        RECT 118.255 190.875 119.465 191.625 ;
        RECT 117.225 190.320 117.500 190.650 ;
        RECT 117.725 190.355 118.065 190.725 ;
        RECT 117.330 190.175 117.500 190.320 ;
        RECT 111.355 189.075 116.700 189.510 ;
        RECT 116.875 189.245 117.145 190.150 ;
        RECT 117.330 190.005 118.005 190.175 ;
        RECT 117.315 189.075 117.645 189.835 ;
        RECT 117.825 189.245 118.005 190.005 ;
        RECT 118.255 190.165 118.775 190.705 ;
        RECT 118.945 190.335 119.465 190.875 ;
        RECT 118.255 189.075 119.465 190.165 ;
        RECT 71.250 188.905 119.550 189.075 ;
        RECT 71.335 187.815 72.545 188.905 ;
        RECT 72.715 188.470 78.060 188.905 ;
        RECT 71.335 187.105 71.855 187.645 ;
        RECT 72.025 187.275 72.545 187.815 ;
        RECT 71.335 186.355 72.545 187.105 ;
        RECT 74.300 186.900 74.640 187.730 ;
        RECT 76.120 187.220 76.470 188.470 ;
        RECT 78.235 187.815 79.905 188.905 ;
        RECT 80.535 187.830 80.875 188.905 ;
        RECT 81.060 188.395 83.110 188.685 ;
        RECT 78.235 187.125 78.985 187.645 ;
        RECT 79.155 187.295 79.905 187.815 ;
        RECT 81.045 187.595 81.285 188.190 ;
        RECT 81.480 188.055 83.110 188.225 ;
        RECT 83.280 188.105 83.560 188.905 ;
        RECT 81.480 187.765 81.800 188.055 ;
        RECT 82.940 187.935 83.110 188.055 ;
        RECT 72.715 186.355 78.060 186.900 ;
        RECT 78.235 186.355 79.905 187.125 ;
        RECT 80.535 187.025 80.875 187.595 ;
        RECT 81.045 187.265 81.700 187.595 ;
        RECT 81.970 187.265 82.710 187.885 ;
        RECT 82.940 187.765 83.600 187.935 ;
        RECT 83.770 187.765 84.045 188.735 ;
        RECT 83.430 187.595 83.600 187.765 ;
        RECT 82.880 187.265 83.260 187.595 ;
        RECT 83.430 187.265 83.705 187.595 ;
        RECT 80.535 186.355 80.875 186.855 ;
        RECT 81.045 186.575 81.290 187.265 ;
        RECT 83.430 187.095 83.600 187.265 ;
        RECT 82.015 186.925 83.600 187.095 ;
        RECT 83.875 187.030 84.045 187.765 ;
        RECT 84.215 187.740 84.505 188.905 ;
        RECT 84.765 188.235 84.935 188.735 ;
        RECT 85.105 188.405 85.435 188.905 ;
        RECT 84.765 188.065 85.430 188.235 ;
        RECT 84.680 187.245 85.030 187.895 ;
        RECT 81.485 186.355 81.815 186.855 ;
        RECT 82.015 186.575 82.185 186.925 ;
        RECT 82.360 186.355 82.690 186.755 ;
        RECT 82.860 186.575 83.030 186.925 ;
        RECT 83.200 186.355 83.580 186.755 ;
        RECT 83.770 186.685 84.045 187.030 ;
        RECT 84.215 186.355 84.505 187.080 ;
        RECT 85.200 187.075 85.430 188.065 ;
        RECT 84.765 186.905 85.430 187.075 ;
        RECT 84.765 186.615 84.935 186.905 ;
        RECT 85.105 186.355 85.435 186.735 ;
        RECT 85.605 186.615 85.790 188.735 ;
        RECT 86.030 188.445 86.295 188.905 ;
        RECT 86.465 188.310 86.715 188.735 ;
        RECT 86.925 188.460 88.030 188.630 ;
        RECT 86.410 188.180 86.715 188.310 ;
        RECT 85.960 186.985 86.240 187.935 ;
        RECT 86.410 187.075 86.580 188.180 ;
        RECT 86.750 187.395 86.990 187.990 ;
        RECT 87.160 187.925 87.690 188.290 ;
        RECT 87.160 187.225 87.330 187.925 ;
        RECT 87.860 187.845 88.030 188.460 ;
        RECT 88.200 188.105 88.370 188.905 ;
        RECT 88.540 188.405 88.790 188.735 ;
        RECT 89.015 188.435 89.900 188.605 ;
        RECT 87.860 187.755 88.370 187.845 ;
        RECT 86.410 186.945 86.635 187.075 ;
        RECT 86.805 187.005 87.330 187.225 ;
        RECT 87.500 187.585 88.370 187.755 ;
        RECT 86.045 186.355 86.295 186.815 ;
        RECT 86.465 186.805 86.635 186.945 ;
        RECT 87.500 186.805 87.670 187.585 ;
        RECT 88.200 187.515 88.370 187.585 ;
        RECT 87.880 187.335 88.080 187.365 ;
        RECT 88.540 187.335 88.710 188.405 ;
        RECT 88.880 187.515 89.070 188.235 ;
        RECT 87.880 187.035 88.710 187.335 ;
        RECT 89.240 187.305 89.560 188.265 ;
        RECT 86.465 186.635 86.800 186.805 ;
        RECT 86.995 186.635 87.670 186.805 ;
        RECT 87.990 186.355 88.360 186.855 ;
        RECT 88.540 186.805 88.710 187.035 ;
        RECT 89.095 186.975 89.560 187.305 ;
        RECT 89.730 187.595 89.900 188.435 ;
        RECT 90.080 188.405 90.395 188.905 ;
        RECT 90.625 188.175 90.965 188.735 ;
        RECT 90.070 187.800 90.965 188.175 ;
        RECT 91.135 187.895 91.305 188.905 ;
        RECT 90.775 187.595 90.965 187.800 ;
        RECT 91.475 187.845 91.805 188.690 ;
        RECT 91.475 187.765 91.865 187.845 ;
        RECT 91.650 187.715 91.865 187.765 ;
        RECT 89.730 187.265 90.605 187.595 ;
        RECT 90.775 187.265 91.525 187.595 ;
        RECT 89.730 186.805 89.900 187.265 ;
        RECT 90.775 187.095 90.975 187.265 ;
        RECT 91.695 187.135 91.865 187.715 ;
        RECT 91.640 187.095 91.865 187.135 ;
        RECT 88.540 186.635 88.945 186.805 ;
        RECT 89.115 186.635 89.900 186.805 ;
        RECT 90.175 186.355 90.385 186.885 ;
        RECT 90.645 186.570 90.975 187.095 ;
        RECT 91.485 187.010 91.865 187.095 ;
        RECT 92.035 187.765 92.420 188.735 ;
        RECT 92.590 188.445 92.915 188.905 ;
        RECT 93.435 188.275 93.715 188.735 ;
        RECT 92.590 188.055 93.715 188.275 ;
        RECT 92.035 187.095 92.315 187.765 ;
        RECT 92.590 187.595 93.040 188.055 ;
        RECT 93.905 187.885 94.305 188.735 ;
        RECT 94.705 188.445 94.975 188.905 ;
        RECT 95.145 188.275 95.430 188.735 ;
        RECT 92.485 187.265 93.040 187.595 ;
        RECT 93.210 187.325 94.305 187.885 ;
        RECT 92.590 187.155 93.040 187.265 ;
        RECT 91.145 186.355 91.315 186.965 ;
        RECT 91.485 186.575 91.815 187.010 ;
        RECT 92.035 186.525 92.420 187.095 ;
        RECT 92.590 186.985 93.715 187.155 ;
        RECT 92.590 186.355 92.915 186.815 ;
        RECT 93.435 186.525 93.715 186.985 ;
        RECT 93.905 186.525 94.305 187.325 ;
        RECT 94.475 188.055 95.430 188.275 ;
        RECT 94.475 187.155 94.685 188.055 ;
        RECT 94.855 187.325 95.545 187.885 ;
        RECT 95.755 187.765 95.985 188.905 ;
        RECT 96.155 187.755 96.485 188.735 ;
        RECT 96.655 187.765 96.865 188.905 ;
        RECT 97.185 188.235 97.355 188.735 ;
        RECT 97.525 188.405 97.855 188.905 ;
        RECT 97.185 188.065 97.850 188.235 ;
        RECT 95.735 187.345 96.065 187.595 ;
        RECT 94.475 186.985 95.430 187.155 ;
        RECT 94.705 186.355 94.975 186.815 ;
        RECT 95.145 186.525 95.430 186.985 ;
        RECT 95.755 186.355 95.985 187.175 ;
        RECT 96.235 187.155 96.485 187.755 ;
        RECT 97.100 187.245 97.450 187.895 ;
        RECT 96.155 186.525 96.485 187.155 ;
        RECT 96.655 186.355 96.865 187.175 ;
        RECT 97.620 187.075 97.850 188.065 ;
        RECT 97.185 186.905 97.850 187.075 ;
        RECT 97.185 186.615 97.355 186.905 ;
        RECT 97.525 186.355 97.855 186.735 ;
        RECT 98.025 186.615 98.210 188.735 ;
        RECT 98.450 188.445 98.715 188.905 ;
        RECT 98.885 188.310 99.135 188.735 ;
        RECT 99.345 188.460 100.450 188.630 ;
        RECT 98.830 188.180 99.135 188.310 ;
        RECT 98.380 186.985 98.660 187.935 ;
        RECT 98.830 187.075 99.000 188.180 ;
        RECT 99.170 187.395 99.410 187.990 ;
        RECT 99.580 187.925 100.110 188.290 ;
        RECT 99.580 187.225 99.750 187.925 ;
        RECT 100.280 187.845 100.450 188.460 ;
        RECT 100.620 188.105 100.790 188.905 ;
        RECT 100.960 188.405 101.210 188.735 ;
        RECT 101.435 188.435 102.320 188.605 ;
        RECT 100.280 187.755 100.790 187.845 ;
        RECT 98.830 186.945 99.055 187.075 ;
        RECT 99.225 187.005 99.750 187.225 ;
        RECT 99.920 187.585 100.790 187.755 ;
        RECT 98.465 186.355 98.715 186.815 ;
        RECT 98.885 186.805 99.055 186.945 ;
        RECT 99.920 186.805 100.090 187.585 ;
        RECT 100.620 187.515 100.790 187.585 ;
        RECT 100.300 187.335 100.500 187.365 ;
        RECT 100.960 187.335 101.130 188.405 ;
        RECT 101.300 187.515 101.490 188.235 ;
        RECT 100.300 187.035 101.130 187.335 ;
        RECT 101.660 187.305 101.980 188.265 ;
        RECT 98.885 186.635 99.220 186.805 ;
        RECT 99.415 186.635 100.090 186.805 ;
        RECT 100.410 186.355 100.780 186.855 ;
        RECT 100.960 186.805 101.130 187.035 ;
        RECT 101.515 186.975 101.980 187.305 ;
        RECT 102.150 187.595 102.320 188.435 ;
        RECT 102.500 188.405 102.815 188.905 ;
        RECT 103.045 188.175 103.385 188.735 ;
        RECT 102.490 187.800 103.385 188.175 ;
        RECT 103.555 187.895 103.725 188.905 ;
        RECT 103.195 187.595 103.385 187.800 ;
        RECT 103.895 187.845 104.225 188.690 ;
        RECT 104.455 188.105 104.895 188.735 ;
        RECT 103.895 187.765 104.285 187.845 ;
        RECT 104.070 187.715 104.285 187.765 ;
        RECT 102.150 187.265 103.025 187.595 ;
        RECT 103.195 187.265 103.945 187.595 ;
        RECT 102.150 186.805 102.320 187.265 ;
        RECT 103.195 187.095 103.395 187.265 ;
        RECT 104.115 187.135 104.285 187.715 ;
        RECT 104.060 187.095 104.285 187.135 ;
        RECT 100.960 186.635 101.365 186.805 ;
        RECT 101.535 186.635 102.320 186.805 ;
        RECT 102.595 186.355 102.805 186.885 ;
        RECT 103.065 186.570 103.395 187.095 ;
        RECT 103.905 187.010 104.285 187.095 ;
        RECT 104.455 187.095 104.765 188.105 ;
        RECT 105.070 188.055 105.385 188.905 ;
        RECT 105.555 188.565 106.985 188.735 ;
        RECT 105.555 187.885 105.725 188.565 ;
        RECT 104.935 187.715 105.725 187.885 ;
        RECT 104.935 187.265 105.105 187.715 ;
        RECT 105.895 187.595 106.095 188.395 ;
        RECT 105.275 187.265 105.665 187.545 ;
        RECT 105.850 187.265 106.095 187.595 ;
        RECT 106.295 187.265 106.545 188.395 ;
        RECT 106.735 187.935 106.985 188.565 ;
        RECT 107.165 188.105 107.495 188.905 ;
        RECT 107.685 187.935 108.015 188.720 ;
        RECT 106.735 187.765 107.505 187.935 ;
        RECT 107.685 187.765 108.365 187.935 ;
        RECT 108.545 187.765 108.875 188.905 ;
        RECT 106.760 187.265 107.165 187.595 ;
        RECT 107.335 187.095 107.505 187.765 ;
        RECT 107.675 187.345 108.025 187.595 ;
        RECT 108.195 187.165 108.365 187.765 ;
        RECT 109.975 187.740 110.265 188.905 ;
        RECT 111.360 187.765 111.615 188.905 ;
        RECT 111.810 188.355 113.005 188.685 ;
        RECT 111.865 187.595 112.035 188.155 ;
        RECT 112.260 187.935 112.680 188.185 ;
        RECT 113.185 188.105 113.465 188.905 ;
        RECT 112.260 187.765 113.505 187.935 ;
        RECT 113.675 187.765 113.945 188.735 ;
        RECT 113.335 187.595 113.505 187.765 ;
        RECT 113.715 187.715 113.945 187.765 ;
        RECT 108.535 187.345 108.885 187.595 ;
        RECT 111.360 187.345 111.695 187.595 ;
        RECT 111.865 187.265 112.605 187.595 ;
        RECT 113.335 187.265 113.565 187.595 ;
        RECT 111.865 187.175 112.115 187.265 ;
        RECT 103.565 186.355 103.735 186.965 ;
        RECT 103.905 186.575 104.235 187.010 ;
        RECT 104.455 186.535 104.895 187.095 ;
        RECT 105.065 186.355 105.515 187.095 ;
        RECT 105.685 186.925 106.845 187.095 ;
        RECT 105.685 186.525 105.855 186.925 ;
        RECT 106.025 186.355 106.445 186.755 ;
        RECT 106.615 186.525 106.845 186.925 ;
        RECT 107.015 186.525 107.505 187.095 ;
        RECT 107.695 186.355 107.935 187.165 ;
        RECT 108.105 186.525 108.435 187.165 ;
        RECT 108.605 186.355 108.875 187.165 ;
        RECT 109.975 186.355 110.265 187.080 ;
        RECT 111.380 187.005 112.115 187.175 ;
        RECT 113.335 187.095 113.505 187.265 ;
        RECT 111.380 186.535 111.690 187.005 ;
        RECT 112.765 186.925 113.505 187.095 ;
        RECT 113.775 187.030 113.945 187.715 ;
        RECT 111.860 186.355 112.595 186.835 ;
        RECT 112.765 186.575 112.935 186.925 ;
        RECT 113.105 186.355 113.485 186.755 ;
        RECT 113.675 186.685 113.945 187.030 ;
        RECT 114.115 187.830 114.385 188.735 ;
        RECT 114.555 188.145 114.885 188.905 ;
        RECT 115.065 187.975 115.235 188.735 ;
        RECT 114.115 187.030 114.285 187.830 ;
        RECT 114.570 187.805 115.235 187.975 ;
        RECT 115.495 187.815 118.085 188.905 ;
        RECT 114.570 187.660 114.740 187.805 ;
        RECT 114.455 187.330 114.740 187.660 ;
        RECT 114.570 187.075 114.740 187.330 ;
        RECT 114.975 187.255 115.305 187.625 ;
        RECT 115.495 187.125 116.705 187.645 ;
        RECT 116.875 187.295 118.085 187.815 ;
        RECT 118.255 187.815 119.465 188.905 ;
        RECT 118.255 187.275 118.775 187.815 ;
        RECT 114.115 186.525 114.375 187.030 ;
        RECT 114.570 186.905 115.235 187.075 ;
        RECT 114.555 186.355 114.885 186.735 ;
        RECT 115.065 186.525 115.235 186.905 ;
        RECT 115.495 186.355 118.085 187.125 ;
        RECT 118.945 187.105 119.465 187.645 ;
        RECT 118.255 186.355 119.465 187.105 ;
        RECT 71.250 186.185 119.550 186.355 ;
        RECT 71.335 185.435 72.545 186.185 ;
        RECT 72.715 185.640 78.060 186.185 ;
        RECT 78.235 185.640 83.580 186.185 ;
        RECT 71.335 184.895 71.855 185.435 ;
        RECT 72.025 184.725 72.545 185.265 ;
        RECT 74.300 184.810 74.640 185.640 ;
        RECT 71.335 183.635 72.545 184.725 ;
        RECT 76.120 184.070 76.470 185.320 ;
        RECT 79.820 184.810 80.160 185.640 ;
        RECT 83.755 185.510 84.030 185.855 ;
        RECT 84.220 185.785 84.595 186.185 ;
        RECT 84.765 185.615 84.935 185.965 ;
        RECT 85.105 185.785 85.435 186.185 ;
        RECT 85.605 185.615 85.865 186.015 ;
        RECT 81.640 184.070 81.990 185.320 ;
        RECT 83.755 184.775 83.925 185.510 ;
        RECT 84.200 185.445 85.865 185.615 ;
        RECT 84.200 185.275 84.370 185.445 ;
        RECT 86.045 185.365 86.375 185.785 ;
        RECT 86.545 185.365 86.805 186.185 ;
        RECT 86.975 185.445 87.235 186.015 ;
        RECT 87.405 185.785 87.790 186.185 ;
        RECT 87.960 185.615 88.215 186.015 ;
        RECT 87.405 185.445 88.215 185.615 ;
        RECT 88.405 185.445 88.650 186.015 ;
        RECT 88.820 185.785 89.205 186.185 ;
        RECT 89.375 185.615 89.630 186.015 ;
        RECT 88.820 185.445 89.630 185.615 ;
        RECT 89.820 185.445 90.245 186.015 ;
        RECT 90.415 185.785 90.800 186.185 ;
        RECT 90.970 185.615 91.405 186.015 ;
        RECT 90.415 185.445 91.405 185.615 ;
        RECT 86.045 185.275 86.295 185.365 ;
        RECT 84.095 184.945 84.370 185.275 ;
        RECT 84.540 184.945 85.365 185.275 ;
        RECT 85.580 184.945 86.295 185.275 ;
        RECT 86.465 184.945 86.800 185.195 ;
        RECT 84.200 184.775 84.370 184.945 ;
        RECT 72.715 183.635 78.060 184.070 ;
        RECT 78.235 183.635 83.580 184.070 ;
        RECT 83.755 183.805 84.030 184.775 ;
        RECT 84.200 184.605 84.860 184.775 ;
        RECT 85.120 184.655 85.365 184.945 ;
        RECT 84.690 184.485 84.860 184.605 ;
        RECT 85.535 184.485 85.865 184.775 ;
        RECT 84.240 183.635 84.520 184.435 ;
        RECT 84.690 184.315 85.865 184.485 ;
        RECT 86.125 184.385 86.295 184.945 ;
        RECT 86.975 184.775 87.160 185.445 ;
        RECT 87.405 185.275 87.755 185.445 ;
        RECT 88.405 185.275 88.575 185.445 ;
        RECT 88.820 185.275 89.170 185.445 ;
        RECT 89.820 185.275 90.170 185.445 ;
        RECT 90.415 185.275 90.750 185.445 ;
        RECT 91.575 185.415 93.245 186.185 ;
        RECT 93.530 185.555 93.815 186.015 ;
        RECT 93.985 185.725 94.255 186.185 ;
        RECT 87.330 184.945 87.755 185.275 ;
        RECT 84.690 183.815 86.305 184.145 ;
        RECT 86.545 183.635 86.805 184.775 ;
        RECT 86.975 183.805 87.235 184.775 ;
        RECT 87.405 184.425 87.755 184.945 ;
        RECT 87.925 184.775 88.575 185.275 ;
        RECT 88.745 184.945 89.170 185.275 ;
        RECT 87.925 184.595 88.650 184.775 ;
        RECT 87.405 184.230 88.215 184.425 ;
        RECT 87.405 183.635 87.790 184.060 ;
        RECT 87.960 183.805 88.215 184.230 ;
        RECT 88.405 183.805 88.650 184.595 ;
        RECT 88.820 184.425 89.170 184.945 ;
        RECT 89.340 184.775 90.170 185.275 ;
        RECT 90.340 184.945 90.750 185.275 ;
        RECT 89.340 184.595 90.245 184.775 ;
        RECT 88.820 184.230 89.650 184.425 ;
        RECT 88.820 183.635 89.205 184.060 ;
        RECT 89.375 183.805 89.650 184.230 ;
        RECT 89.820 183.805 90.245 184.595 ;
        RECT 90.415 184.400 90.750 184.945 ;
        RECT 90.920 184.570 91.405 185.275 ;
        RECT 91.575 184.895 92.325 185.415 ;
        RECT 93.530 185.385 94.485 185.555 ;
        RECT 92.495 184.725 93.245 185.245 ;
        RECT 90.415 184.230 91.405 184.400 ;
        RECT 90.415 183.635 90.800 184.060 ;
        RECT 90.970 183.805 91.405 184.230 ;
        RECT 91.575 183.635 93.245 184.725 ;
        RECT 93.415 184.655 94.105 185.215 ;
        RECT 94.275 184.485 94.485 185.385 ;
        RECT 93.530 184.265 94.485 184.485 ;
        RECT 94.655 185.215 95.055 186.015 ;
        RECT 95.245 185.555 95.525 186.015 ;
        RECT 96.045 185.725 96.370 186.185 ;
        RECT 95.245 185.385 96.370 185.555 ;
        RECT 96.540 185.445 96.925 186.015 ;
        RECT 97.095 185.460 97.385 186.185 ;
        RECT 95.920 185.275 96.370 185.385 ;
        RECT 94.655 184.655 95.750 185.215 ;
        RECT 95.920 184.945 96.475 185.275 ;
        RECT 93.530 183.805 93.815 184.265 ;
        RECT 93.985 183.635 94.255 184.095 ;
        RECT 94.655 183.805 95.055 184.655 ;
        RECT 95.920 184.485 96.370 184.945 ;
        RECT 96.645 184.775 96.925 185.445 ;
        RECT 98.475 185.445 98.815 186.015 ;
        RECT 99.010 185.520 99.180 186.185 ;
        RECT 99.460 185.845 99.680 185.890 ;
        RECT 99.455 185.675 99.680 185.845 ;
        RECT 99.850 185.705 100.295 185.875 ;
        RECT 99.460 185.535 99.680 185.675 ;
        RECT 95.245 184.265 96.370 184.485 ;
        RECT 95.245 183.805 95.525 184.265 ;
        RECT 96.045 183.635 96.370 184.095 ;
        RECT 96.540 183.805 96.925 184.775 ;
        RECT 97.095 183.635 97.385 184.800 ;
        RECT 98.475 184.475 98.650 185.445 ;
        RECT 99.460 185.365 99.955 185.535 ;
        RECT 98.820 184.825 98.990 185.275 ;
        RECT 99.160 184.995 99.610 185.195 ;
        RECT 99.780 185.170 99.955 185.365 ;
        RECT 100.125 184.915 100.295 185.705 ;
        RECT 100.465 185.580 100.715 185.950 ;
        RECT 100.545 185.195 100.715 185.580 ;
        RECT 100.885 185.545 101.135 185.950 ;
        RECT 101.305 185.715 101.475 186.185 ;
        RECT 101.645 185.545 101.985 185.950 ;
        RECT 100.885 185.365 101.985 185.545 ;
        RECT 102.170 185.615 102.425 185.965 ;
        RECT 102.595 185.785 102.925 186.185 ;
        RECT 103.095 185.615 103.265 185.965 ;
        RECT 103.435 185.785 103.815 186.185 ;
        RECT 102.170 185.445 103.835 185.615 ;
        RECT 104.005 185.510 104.280 185.855 ;
        RECT 103.665 185.275 103.835 185.445 ;
        RECT 100.545 185.025 100.740 185.195 ;
        RECT 98.820 184.655 99.215 184.825 ;
        RECT 100.125 184.775 100.400 184.915 ;
        RECT 98.475 183.805 98.735 184.475 ;
        RECT 99.045 184.385 99.215 184.655 ;
        RECT 99.385 184.555 100.400 184.775 ;
        RECT 100.570 184.775 100.740 185.025 ;
        RECT 100.910 184.945 101.470 185.195 ;
        RECT 100.570 184.385 101.125 184.775 ;
        RECT 99.045 184.215 101.125 184.385 ;
        RECT 98.905 183.635 99.235 184.035 ;
        RECT 100.105 183.635 100.505 184.035 ;
        RECT 100.795 183.980 101.125 184.215 ;
        RECT 101.295 183.845 101.470 184.945 ;
        RECT 101.640 184.625 101.985 185.195 ;
        RECT 102.155 184.945 102.500 185.275 ;
        RECT 102.670 184.945 103.495 185.275 ;
        RECT 103.665 184.945 103.940 185.275 ;
        RECT 102.175 184.485 102.500 184.775 ;
        RECT 102.670 184.655 102.865 184.945 ;
        RECT 103.665 184.775 103.835 184.945 ;
        RECT 104.110 184.775 104.280 185.510 ;
        RECT 104.455 185.415 106.125 186.185 ;
        RECT 106.295 185.510 106.555 186.015 ;
        RECT 106.735 185.805 107.065 186.185 ;
        RECT 107.245 185.635 107.415 186.015 ;
        RECT 104.455 184.895 105.205 185.415 ;
        RECT 103.175 184.605 103.835 184.775 ;
        RECT 103.175 184.485 103.345 184.605 ;
        RECT 101.640 183.635 101.985 184.455 ;
        RECT 102.175 184.315 103.345 184.485 ;
        RECT 102.155 183.855 103.345 184.145 ;
        RECT 103.515 183.635 103.795 184.435 ;
        RECT 104.005 183.805 104.280 184.775 ;
        RECT 105.375 184.725 106.125 185.245 ;
        RECT 104.455 183.635 106.125 184.725 ;
        RECT 106.295 184.710 106.465 185.510 ;
        RECT 106.750 185.465 107.415 185.635 ;
        RECT 107.675 185.510 107.935 186.015 ;
        RECT 108.115 185.805 108.445 186.185 ;
        RECT 108.625 185.635 108.795 186.015 ;
        RECT 106.750 185.210 106.920 185.465 ;
        RECT 106.635 184.880 106.920 185.210 ;
        RECT 107.155 184.915 107.485 185.285 ;
        RECT 106.750 184.735 106.920 184.880 ;
        RECT 106.295 183.805 106.565 184.710 ;
        RECT 106.750 184.565 107.415 184.735 ;
        RECT 106.735 183.635 107.065 184.395 ;
        RECT 107.245 183.805 107.415 184.565 ;
        RECT 107.675 184.710 107.845 185.510 ;
        RECT 108.130 185.465 108.795 185.635 ;
        RECT 108.130 185.210 108.300 185.465 ;
        RECT 109.055 185.415 110.725 186.185 ;
        RECT 110.985 185.635 111.155 185.925 ;
        RECT 111.325 185.805 111.655 186.185 ;
        RECT 110.985 185.465 111.650 185.635 ;
        RECT 108.015 184.880 108.300 185.210 ;
        RECT 108.535 184.915 108.865 185.285 ;
        RECT 109.055 184.895 109.805 185.415 ;
        RECT 108.130 184.735 108.300 184.880 ;
        RECT 107.675 183.805 107.945 184.710 ;
        RECT 108.130 184.565 108.795 184.735 ;
        RECT 109.975 184.725 110.725 185.245 ;
        RECT 108.115 183.635 108.445 184.395 ;
        RECT 108.625 183.805 108.795 184.565 ;
        RECT 109.055 183.635 110.725 184.725 ;
        RECT 110.900 184.645 111.250 185.295 ;
        RECT 111.420 184.475 111.650 185.465 ;
        RECT 110.985 184.305 111.650 184.475 ;
        RECT 110.985 183.805 111.155 184.305 ;
        RECT 111.325 183.635 111.655 184.135 ;
        RECT 111.825 183.805 112.010 185.925 ;
        RECT 112.265 185.725 112.515 186.185 ;
        RECT 112.685 185.735 113.020 185.905 ;
        RECT 113.215 185.735 113.890 185.905 ;
        RECT 112.685 185.595 112.855 185.735 ;
        RECT 112.180 184.605 112.460 185.555 ;
        RECT 112.630 185.465 112.855 185.595 ;
        RECT 112.630 184.360 112.800 185.465 ;
        RECT 113.025 185.315 113.550 185.535 ;
        RECT 112.970 184.550 113.210 185.145 ;
        RECT 113.380 184.615 113.550 185.315 ;
        RECT 113.720 184.955 113.890 185.735 ;
        RECT 114.210 185.685 114.580 186.185 ;
        RECT 114.760 185.735 115.165 185.905 ;
        RECT 115.335 185.735 116.120 185.905 ;
        RECT 114.760 185.505 114.930 185.735 ;
        RECT 114.100 185.205 114.930 185.505 ;
        RECT 115.315 185.235 115.780 185.565 ;
        RECT 114.100 185.175 114.300 185.205 ;
        RECT 114.420 184.955 114.590 185.025 ;
        RECT 113.720 184.785 114.590 184.955 ;
        RECT 114.080 184.695 114.590 184.785 ;
        RECT 112.630 184.230 112.935 184.360 ;
        RECT 113.380 184.250 113.910 184.615 ;
        RECT 112.250 183.635 112.515 184.095 ;
        RECT 112.685 183.805 112.935 184.230 ;
        RECT 114.080 184.080 114.250 184.695 ;
        RECT 113.145 183.910 114.250 184.080 ;
        RECT 114.420 183.635 114.590 184.435 ;
        RECT 114.760 184.135 114.930 185.205 ;
        RECT 115.100 184.305 115.290 185.025 ;
        RECT 115.460 184.275 115.780 185.235 ;
        RECT 115.950 185.275 116.120 185.735 ;
        RECT 116.395 185.655 116.605 186.185 ;
        RECT 116.865 185.445 117.195 185.970 ;
        RECT 117.365 185.575 117.535 186.185 ;
        RECT 117.705 185.530 118.035 185.965 ;
        RECT 117.705 185.445 118.085 185.530 ;
        RECT 116.995 185.275 117.195 185.445 ;
        RECT 117.860 185.405 118.085 185.445 ;
        RECT 118.255 185.435 119.465 186.185 ;
        RECT 115.950 184.945 116.825 185.275 ;
        RECT 116.995 184.945 117.745 185.275 ;
        RECT 114.760 183.805 115.010 184.135 ;
        RECT 115.950 184.105 116.120 184.945 ;
        RECT 116.995 184.740 117.185 184.945 ;
        RECT 117.915 184.825 118.085 185.405 ;
        RECT 117.870 184.775 118.085 184.825 ;
        RECT 116.290 184.365 117.185 184.740 ;
        RECT 117.695 184.695 118.085 184.775 ;
        RECT 118.255 184.725 118.775 185.265 ;
        RECT 118.945 184.895 119.465 185.435 ;
        RECT 115.235 183.935 116.120 184.105 ;
        RECT 116.300 183.635 116.615 184.135 ;
        RECT 116.845 183.805 117.185 184.365 ;
        RECT 117.355 183.635 117.525 184.645 ;
        RECT 117.695 183.850 118.025 184.695 ;
        RECT 118.255 183.635 119.465 184.725 ;
        RECT 71.250 183.465 119.550 183.635 ;
        RECT 71.335 182.375 72.545 183.465 ;
        RECT 72.715 183.030 78.060 183.465 ;
        RECT 78.235 183.030 83.580 183.465 ;
        RECT 71.335 181.665 71.855 182.205 ;
        RECT 72.025 181.835 72.545 182.375 ;
        RECT 71.335 180.915 72.545 181.665 ;
        RECT 74.300 181.460 74.640 182.290 ;
        RECT 76.120 181.780 76.470 183.030 ;
        RECT 79.820 181.460 80.160 182.290 ;
        RECT 81.640 181.780 81.990 183.030 ;
        RECT 84.215 182.300 84.505 183.465 ;
        RECT 84.675 182.375 86.345 183.465 ;
        RECT 87.090 182.835 87.375 183.295 ;
        RECT 87.545 183.005 87.815 183.465 ;
        RECT 87.090 182.615 88.045 182.835 ;
        RECT 84.675 181.685 85.425 182.205 ;
        RECT 85.595 181.855 86.345 182.375 ;
        RECT 86.975 181.885 87.665 182.445 ;
        RECT 87.835 181.715 88.045 182.615 ;
        RECT 72.715 180.915 78.060 181.460 ;
        RECT 78.235 180.915 83.580 181.460 ;
        RECT 84.215 180.915 84.505 181.640 ;
        RECT 84.675 180.915 86.345 181.685 ;
        RECT 87.090 181.545 88.045 181.715 ;
        RECT 88.215 182.445 88.615 183.295 ;
        RECT 88.805 182.835 89.085 183.295 ;
        RECT 89.605 183.005 89.930 183.465 ;
        RECT 88.805 182.615 89.930 182.835 ;
        RECT 88.215 181.885 89.310 182.445 ;
        RECT 89.480 182.155 89.930 182.615 ;
        RECT 90.100 182.325 90.485 183.295 ;
        RECT 90.655 182.375 92.325 183.465 ;
        RECT 87.090 181.085 87.375 181.545 ;
        RECT 87.545 180.915 87.815 181.375 ;
        RECT 88.215 181.085 88.615 181.885 ;
        RECT 89.480 181.825 90.035 182.155 ;
        RECT 89.480 181.715 89.930 181.825 ;
        RECT 88.805 181.545 89.930 181.715 ;
        RECT 90.205 181.655 90.485 182.325 ;
        RECT 88.805 181.085 89.085 181.545 ;
        RECT 89.605 180.915 89.930 181.375 ;
        RECT 90.100 181.085 90.485 181.655 ;
        RECT 90.655 181.685 91.405 182.205 ;
        RECT 91.575 181.855 92.325 182.375 ;
        RECT 92.500 182.325 92.755 183.465 ;
        RECT 92.950 182.915 94.145 183.245 ;
        RECT 93.005 182.155 93.175 182.715 ;
        RECT 93.400 182.495 93.820 182.745 ;
        RECT 94.325 182.665 94.605 183.465 ;
        RECT 93.400 182.325 94.645 182.495 ;
        RECT 94.815 182.325 95.085 183.295 ;
        RECT 95.715 182.325 95.975 183.465 ;
        RECT 96.145 182.495 96.475 183.295 ;
        RECT 96.645 182.665 96.815 183.465 ;
        RECT 96.985 182.495 97.315 183.295 ;
        RECT 97.485 182.665 97.740 183.465 ;
        RECT 98.015 183.030 103.360 183.465 ;
        RECT 96.145 182.325 97.845 182.495 ;
        RECT 94.475 182.155 94.645 182.325 ;
        RECT 92.500 181.905 92.835 182.155 ;
        RECT 93.005 181.825 93.745 182.155 ;
        RECT 94.475 181.825 94.705 182.155 ;
        RECT 93.005 181.735 93.255 181.825 ;
        RECT 90.655 180.915 92.325 181.685 ;
        RECT 92.520 181.565 93.255 181.735 ;
        RECT 94.475 181.655 94.645 181.825 ;
        RECT 92.520 181.095 92.830 181.565 ;
        RECT 93.905 181.485 94.645 181.655 ;
        RECT 94.915 181.590 95.085 182.325 ;
        RECT 95.715 181.905 96.475 182.155 ;
        RECT 96.645 181.905 97.395 182.155 ;
        RECT 97.565 181.735 97.845 182.325 ;
        RECT 93.000 180.915 93.735 181.395 ;
        RECT 93.905 181.135 94.075 181.485 ;
        RECT 94.245 180.915 94.625 181.315 ;
        RECT 94.815 181.245 95.085 181.590 ;
        RECT 95.715 181.545 96.815 181.715 ;
        RECT 95.715 181.085 96.055 181.545 ;
        RECT 96.225 180.915 96.395 181.375 ;
        RECT 96.565 181.295 96.815 181.545 ;
        RECT 96.985 181.485 97.845 181.735 ;
        RECT 99.600 181.460 99.940 182.290 ;
        RECT 101.420 181.780 101.770 183.030 ;
        RECT 104.100 183.005 104.270 183.465 ;
        RECT 104.440 182.835 104.770 183.295 ;
        RECT 103.995 182.665 104.770 182.835 ;
        RECT 104.940 182.665 105.110 183.465 ;
        RECT 103.995 181.655 104.425 182.665 ;
        RECT 105.695 182.495 106.055 182.670 ;
        RECT 104.595 182.325 106.055 182.495 ;
        RECT 106.295 182.375 109.805 183.465 ;
        RECT 104.595 181.825 104.765 182.325 ;
        RECT 103.995 181.485 104.690 181.655 ;
        RECT 104.935 181.595 105.345 182.155 ;
        RECT 97.405 181.295 97.735 181.315 ;
        RECT 96.565 181.085 97.735 181.295 ;
        RECT 98.015 180.915 103.360 181.460 ;
        RECT 104.020 180.915 104.350 181.315 ;
        RECT 104.520 181.215 104.690 181.485 ;
        RECT 105.515 181.425 105.695 182.325 ;
        RECT 105.865 181.765 106.060 182.155 ;
        RECT 105.865 181.595 106.065 181.765 ;
        RECT 106.295 181.685 107.945 182.205 ;
        RECT 108.115 181.855 109.805 182.375 ;
        RECT 109.975 182.300 110.265 183.465 ;
        RECT 110.435 182.375 113.025 183.465 ;
        RECT 110.435 181.685 111.645 182.205 ;
        RECT 111.815 181.855 113.025 182.375 ;
        RECT 113.255 182.325 113.465 183.465 ;
        RECT 113.635 182.315 113.965 183.295 ;
        RECT 114.135 182.325 114.365 183.465 ;
        RECT 114.575 182.325 114.960 183.295 ;
        RECT 115.130 183.005 115.455 183.465 ;
        RECT 115.975 182.835 116.255 183.295 ;
        RECT 115.130 182.615 116.255 182.835 ;
        RECT 104.860 180.915 105.175 181.425 ;
        RECT 105.405 181.085 105.695 181.425 ;
        RECT 105.865 180.915 106.105 181.425 ;
        RECT 106.295 180.915 109.805 181.685 ;
        RECT 109.975 180.915 110.265 181.640 ;
        RECT 110.435 180.915 113.025 181.685 ;
        RECT 113.255 180.915 113.465 181.735 ;
        RECT 113.635 181.715 113.885 182.315 ;
        RECT 114.055 181.905 114.385 182.155 ;
        RECT 113.635 181.085 113.965 181.715 ;
        RECT 114.135 180.915 114.365 181.735 ;
        RECT 114.575 181.655 114.855 182.325 ;
        RECT 115.130 182.155 115.580 182.615 ;
        RECT 116.445 182.445 116.845 183.295 ;
        RECT 117.245 183.005 117.515 183.465 ;
        RECT 117.685 182.835 117.970 183.295 ;
        RECT 115.025 181.825 115.580 182.155 ;
        RECT 115.750 181.885 116.845 182.445 ;
        RECT 115.130 181.715 115.580 181.825 ;
        RECT 114.575 181.085 114.960 181.655 ;
        RECT 115.130 181.545 116.255 181.715 ;
        RECT 115.130 180.915 115.455 181.375 ;
        RECT 115.975 181.085 116.255 181.545 ;
        RECT 116.445 181.085 116.845 181.885 ;
        RECT 117.015 182.615 117.970 182.835 ;
        RECT 117.015 181.715 117.225 182.615 ;
        RECT 117.395 181.885 118.085 182.445 ;
        RECT 118.255 182.375 119.465 183.465 ;
        RECT 118.255 181.835 118.775 182.375 ;
        RECT 117.015 181.545 117.970 181.715 ;
        RECT 118.945 181.665 119.465 182.205 ;
        RECT 117.245 180.915 117.515 181.375 ;
        RECT 117.685 181.085 117.970 181.545 ;
        RECT 118.255 180.915 119.465 181.665 ;
        RECT 71.250 180.745 119.550 180.915 ;
        RECT 71.335 179.995 72.545 180.745 ;
        RECT 73.640 180.195 73.895 180.485 ;
        RECT 74.065 180.365 74.395 180.745 ;
        RECT 73.640 180.025 74.390 180.195 ;
        RECT 71.335 179.455 71.855 179.995 ;
        RECT 72.025 179.285 72.545 179.825 ;
        RECT 71.335 178.195 72.545 179.285 ;
        RECT 73.640 179.205 73.990 179.855 ;
        RECT 74.160 179.035 74.390 180.025 ;
        RECT 73.640 178.865 74.390 179.035 ;
        RECT 73.640 178.365 73.895 178.865 ;
        RECT 74.065 178.195 74.395 178.695 ;
        RECT 74.565 178.365 74.735 180.485 ;
        RECT 75.095 180.385 75.425 180.745 ;
        RECT 75.595 180.355 76.090 180.525 ;
        RECT 76.295 180.355 77.150 180.525 ;
        RECT 74.965 179.165 75.425 180.215 ;
        RECT 74.905 178.380 75.230 179.165 ;
        RECT 75.595 178.995 75.765 180.355 ;
        RECT 75.935 179.445 76.285 180.065 ;
        RECT 76.455 179.845 76.810 180.065 ;
        RECT 76.455 179.255 76.625 179.845 ;
        RECT 76.980 179.645 77.150 180.355 ;
        RECT 78.025 180.285 78.355 180.745 ;
        RECT 78.565 180.385 78.915 180.555 ;
        RECT 77.355 179.815 78.145 180.065 ;
        RECT 78.565 179.995 78.825 180.385 ;
        RECT 79.135 180.295 80.085 180.575 ;
        RECT 80.255 180.305 80.445 180.745 ;
        RECT 80.615 180.365 81.685 180.535 ;
        RECT 78.315 179.645 78.485 179.825 ;
        RECT 75.595 178.825 75.990 178.995 ;
        RECT 76.160 178.865 76.625 179.255 ;
        RECT 76.795 179.475 78.485 179.645 ;
        RECT 75.820 178.695 75.990 178.825 ;
        RECT 76.795 178.695 76.965 179.475 ;
        RECT 78.655 179.305 78.825 179.995 ;
        RECT 77.325 179.135 78.825 179.305 ;
        RECT 79.015 179.335 79.225 180.125 ;
        RECT 79.395 179.505 79.745 180.125 ;
        RECT 79.915 179.515 80.085 180.295 ;
        RECT 80.615 180.135 80.785 180.365 ;
        RECT 80.255 179.965 80.785 180.135 ;
        RECT 80.255 179.685 80.475 179.965 ;
        RECT 80.955 179.795 81.195 180.195 ;
        RECT 79.915 179.345 80.320 179.515 ;
        RECT 80.655 179.425 81.195 179.795 ;
        RECT 81.365 180.010 81.685 180.365 ;
        RECT 81.930 180.285 82.235 180.745 ;
        RECT 82.405 180.035 82.660 180.565 ;
        RECT 81.365 179.835 81.690 180.010 ;
        RECT 81.365 179.535 82.280 179.835 ;
        RECT 81.540 179.505 82.280 179.535 ;
        RECT 79.015 179.175 79.690 179.335 ;
        RECT 80.150 179.255 80.320 179.345 ;
        RECT 79.015 179.165 79.980 179.175 ;
        RECT 78.655 178.995 78.825 179.135 ;
        RECT 75.400 178.195 75.650 178.655 ;
        RECT 75.820 178.365 76.070 178.695 ;
        RECT 76.285 178.365 76.965 178.695 ;
        RECT 77.135 178.795 78.210 178.965 ;
        RECT 78.655 178.825 79.215 178.995 ;
        RECT 79.520 178.875 79.980 179.165 ;
        RECT 80.150 179.085 81.370 179.255 ;
        RECT 77.135 178.455 77.305 178.795 ;
        RECT 77.540 178.195 77.870 178.625 ;
        RECT 78.040 178.455 78.210 178.795 ;
        RECT 78.505 178.195 78.875 178.655 ;
        RECT 79.045 178.365 79.215 178.825 ;
        RECT 80.150 178.705 80.320 179.085 ;
        RECT 81.540 178.915 81.710 179.505 ;
        RECT 82.450 179.385 82.660 180.035 ;
        RECT 82.835 179.975 84.505 180.745 ;
        RECT 85.135 180.070 85.395 180.575 ;
        RECT 85.575 180.365 85.905 180.745 ;
        RECT 86.085 180.195 86.255 180.575 ;
        RECT 86.515 180.200 91.860 180.745 ;
        RECT 82.835 179.455 83.585 179.975 ;
        RECT 79.450 178.365 80.320 178.705 ;
        RECT 80.910 178.745 81.710 178.915 ;
        RECT 80.490 178.195 80.740 178.655 ;
        RECT 80.910 178.455 81.080 178.745 ;
        RECT 81.260 178.195 81.590 178.575 ;
        RECT 81.930 178.195 82.235 179.335 ;
        RECT 82.405 178.505 82.660 179.385 ;
        RECT 83.755 179.285 84.505 179.805 ;
        RECT 82.835 178.195 84.505 179.285 ;
        RECT 85.135 179.270 85.315 180.070 ;
        RECT 85.590 180.025 86.255 180.195 ;
        RECT 85.590 179.770 85.760 180.025 ;
        RECT 85.485 179.440 85.760 179.770 ;
        RECT 85.985 179.475 86.325 179.845 ;
        RECT 85.590 179.295 85.760 179.440 ;
        RECT 88.100 179.370 88.440 180.200 ;
        RECT 92.035 179.975 95.545 180.745 ;
        RECT 95.715 179.995 96.925 180.745 ;
        RECT 97.095 180.020 97.385 180.745 ;
        RECT 97.590 180.005 98.205 180.575 ;
        RECT 98.375 180.235 98.590 180.745 ;
        RECT 98.820 180.235 99.100 180.565 ;
        RECT 99.280 180.235 99.520 180.745 ;
        RECT 85.135 178.365 85.405 179.270 ;
        RECT 85.590 179.125 86.265 179.295 ;
        RECT 85.575 178.195 85.905 178.955 ;
        RECT 86.085 178.365 86.265 179.125 ;
        RECT 89.920 178.630 90.270 179.880 ;
        RECT 92.035 179.455 93.685 179.975 ;
        RECT 93.855 179.285 95.545 179.805 ;
        RECT 95.715 179.455 96.235 179.995 ;
        RECT 96.405 179.285 96.925 179.825 ;
        RECT 86.515 178.195 91.860 178.630 ;
        RECT 92.035 178.195 95.545 179.285 ;
        RECT 95.715 178.195 96.925 179.285 ;
        RECT 97.095 178.195 97.385 179.360 ;
        RECT 97.590 178.985 97.905 180.005 ;
        RECT 98.075 179.335 98.245 179.835 ;
        RECT 98.495 179.505 98.760 180.065 ;
        RECT 98.930 179.335 99.100 180.235 ;
        RECT 99.270 179.505 99.625 180.065 ;
        RECT 99.855 179.995 101.065 180.745 ;
        RECT 99.855 179.455 100.375 179.995 ;
        RECT 98.075 179.165 99.500 179.335 ;
        RECT 100.545 179.285 101.065 179.825 ;
        RECT 97.590 178.365 98.125 178.985 ;
        RECT 98.295 178.195 98.625 178.995 ;
        RECT 99.110 178.990 99.500 179.165 ;
        RECT 99.855 178.195 101.065 179.285 ;
        RECT 101.245 178.375 101.505 180.565 ;
        RECT 101.765 180.375 102.435 180.745 ;
        RECT 102.615 180.195 102.925 180.565 ;
        RECT 101.695 179.995 102.925 180.195 ;
        RECT 101.695 179.325 101.985 179.995 ;
        RECT 103.105 179.815 103.335 180.455 ;
        RECT 103.515 180.015 103.805 180.745 ;
        RECT 103.995 179.995 105.205 180.745 ;
        RECT 105.465 180.195 105.635 180.485 ;
        RECT 105.805 180.365 106.135 180.745 ;
        RECT 105.465 180.025 106.130 180.195 ;
        RECT 102.165 179.505 102.630 179.815 ;
        RECT 102.810 179.505 103.335 179.815 ;
        RECT 103.515 179.505 103.815 179.835 ;
        RECT 103.995 179.455 104.515 179.995 ;
        RECT 101.695 179.105 102.465 179.325 ;
        RECT 101.675 178.195 102.015 178.925 ;
        RECT 102.195 178.375 102.465 179.105 ;
        RECT 102.645 179.085 103.805 179.325 ;
        RECT 104.685 179.285 105.205 179.825 ;
        RECT 102.645 178.375 102.875 179.085 ;
        RECT 103.045 178.195 103.375 178.905 ;
        RECT 103.545 178.375 103.805 179.085 ;
        RECT 103.995 178.195 105.205 179.285 ;
        RECT 105.380 179.205 105.730 179.855 ;
        RECT 105.900 179.035 106.130 180.025 ;
        RECT 105.465 178.865 106.130 179.035 ;
        RECT 105.465 178.365 105.635 178.865 ;
        RECT 105.805 178.195 106.135 178.695 ;
        RECT 106.305 178.365 106.490 180.485 ;
        RECT 106.745 180.285 106.995 180.745 ;
        RECT 107.165 180.295 107.500 180.465 ;
        RECT 107.695 180.295 108.370 180.465 ;
        RECT 107.165 180.155 107.335 180.295 ;
        RECT 106.660 179.165 106.940 180.115 ;
        RECT 107.110 180.025 107.335 180.155 ;
        RECT 107.110 178.920 107.280 180.025 ;
        RECT 107.505 179.875 108.030 180.095 ;
        RECT 107.450 179.110 107.690 179.705 ;
        RECT 107.860 179.175 108.030 179.875 ;
        RECT 108.200 179.515 108.370 180.295 ;
        RECT 108.690 180.245 109.060 180.745 ;
        RECT 109.240 180.295 109.645 180.465 ;
        RECT 109.815 180.295 110.600 180.465 ;
        RECT 109.240 180.065 109.410 180.295 ;
        RECT 108.580 179.765 109.410 180.065 ;
        RECT 109.795 179.795 110.260 180.125 ;
        RECT 108.580 179.735 108.780 179.765 ;
        RECT 108.900 179.515 109.070 179.585 ;
        RECT 108.200 179.345 109.070 179.515 ;
        RECT 108.560 179.255 109.070 179.345 ;
        RECT 107.110 178.790 107.415 178.920 ;
        RECT 107.860 178.810 108.390 179.175 ;
        RECT 106.730 178.195 106.995 178.655 ;
        RECT 107.165 178.365 107.415 178.790 ;
        RECT 108.560 178.640 108.730 179.255 ;
        RECT 107.625 178.470 108.730 178.640 ;
        RECT 108.900 178.195 109.070 178.995 ;
        RECT 109.240 178.695 109.410 179.765 ;
        RECT 109.580 178.865 109.770 179.585 ;
        RECT 109.940 178.835 110.260 179.795 ;
        RECT 110.430 179.835 110.600 180.295 ;
        RECT 110.875 180.215 111.085 180.745 ;
        RECT 111.345 180.005 111.675 180.530 ;
        RECT 111.845 180.135 112.015 180.745 ;
        RECT 112.185 180.090 112.515 180.525 ;
        RECT 112.735 180.200 118.080 180.745 ;
        RECT 112.185 180.005 112.565 180.090 ;
        RECT 111.475 179.835 111.675 180.005 ;
        RECT 112.340 179.965 112.565 180.005 ;
        RECT 110.430 179.505 111.305 179.835 ;
        RECT 111.475 179.505 112.225 179.835 ;
        RECT 109.240 178.365 109.490 178.695 ;
        RECT 110.430 178.665 110.600 179.505 ;
        RECT 111.475 179.300 111.665 179.505 ;
        RECT 112.395 179.385 112.565 179.965 ;
        RECT 112.350 179.335 112.565 179.385 ;
        RECT 114.320 179.370 114.660 180.200 ;
        RECT 118.255 179.995 119.465 180.745 ;
        RECT 110.770 178.925 111.665 179.300 ;
        RECT 112.175 179.255 112.565 179.335 ;
        RECT 109.715 178.495 110.600 178.665 ;
        RECT 110.780 178.195 111.095 178.695 ;
        RECT 111.325 178.365 111.665 178.925 ;
        RECT 111.835 178.195 112.005 179.205 ;
        RECT 112.175 178.410 112.505 179.255 ;
        RECT 116.140 178.630 116.490 179.880 ;
        RECT 118.255 179.285 118.775 179.825 ;
        RECT 118.945 179.455 119.465 179.995 ;
        RECT 112.735 178.195 118.080 178.630 ;
        RECT 118.255 178.195 119.465 179.285 ;
        RECT 71.250 178.025 119.550 178.195 ;
        RECT 71.335 176.935 72.545 178.025 ;
        RECT 71.335 176.225 71.855 176.765 ;
        RECT 72.025 176.395 72.545 176.935 ;
        RECT 73.635 176.925 73.955 177.855 ;
        RECT 74.135 177.345 74.535 177.855 ;
        RECT 74.705 177.515 74.875 178.025 ;
        RECT 75.045 177.345 75.375 177.855 ;
        RECT 74.135 177.175 75.375 177.345 ;
        RECT 75.545 177.175 75.715 178.025 ;
        RECT 76.305 177.175 76.685 177.855 ;
        RECT 73.635 176.755 74.265 176.925 ;
        RECT 71.335 175.475 72.545 176.225 ;
        RECT 73.635 175.475 73.925 176.310 ;
        RECT 74.095 175.875 74.265 176.755 ;
        RECT 75.040 176.835 76.345 177.005 ;
        RECT 74.435 176.215 74.665 176.715 ;
        RECT 75.040 176.635 75.210 176.835 ;
        RECT 74.835 176.465 75.210 176.635 ;
        RECT 75.380 176.465 75.930 176.665 ;
        RECT 76.100 176.385 76.345 176.835 ;
        RECT 76.515 176.215 76.685 177.175 ;
        RECT 76.855 176.935 80.365 178.025 ;
        RECT 74.435 176.045 76.685 176.215 ;
        RECT 76.855 176.245 78.505 176.765 ;
        RECT 78.675 176.415 80.365 176.935 ;
        RECT 80.995 176.925 81.315 177.855 ;
        RECT 81.495 177.345 81.895 177.855 ;
        RECT 82.065 177.515 82.235 178.025 ;
        RECT 82.405 177.345 82.735 177.855 ;
        RECT 81.495 177.175 82.735 177.345 ;
        RECT 82.905 177.175 83.075 178.025 ;
        RECT 83.665 177.175 84.045 177.855 ;
        RECT 80.995 176.755 81.625 176.925 ;
        RECT 74.095 175.705 75.050 175.875 ;
        RECT 75.465 175.475 75.795 175.865 ;
        RECT 75.965 175.725 76.135 176.045 ;
        RECT 76.305 175.475 76.635 175.865 ;
        RECT 76.855 175.475 80.365 176.245 ;
        RECT 80.995 175.475 81.285 176.310 ;
        RECT 81.455 175.875 81.625 176.755 ;
        RECT 82.400 176.835 83.705 177.005 ;
        RECT 81.795 176.215 82.025 176.715 ;
        RECT 82.400 176.635 82.570 176.835 ;
        RECT 82.195 176.465 82.570 176.635 ;
        RECT 82.740 176.465 83.290 176.665 ;
        RECT 83.460 176.385 83.705 176.835 ;
        RECT 83.875 176.215 84.045 177.175 ;
        RECT 84.215 176.860 84.505 178.025 ;
        RECT 84.675 177.590 90.020 178.025 ;
        RECT 81.795 176.045 84.045 176.215 ;
        RECT 81.455 175.705 82.410 175.875 ;
        RECT 82.825 175.475 83.155 175.865 ;
        RECT 83.325 175.725 83.495 176.045 ;
        RECT 83.665 175.475 83.995 175.865 ;
        RECT 84.215 175.475 84.505 176.200 ;
        RECT 86.260 176.020 86.600 176.850 ;
        RECT 88.080 176.340 88.430 177.590 ;
        RECT 90.195 176.935 91.865 178.025 ;
        RECT 92.045 177.215 92.340 178.025 ;
        RECT 90.195 176.245 90.945 176.765 ;
        RECT 91.115 176.415 91.865 176.935 ;
        RECT 92.520 176.715 92.765 177.855 ;
        RECT 92.940 177.215 93.200 178.025 ;
        RECT 93.800 178.020 100.075 178.025 ;
        RECT 93.380 176.715 93.630 177.850 ;
        RECT 93.800 177.225 94.060 178.020 ;
        RECT 94.230 177.125 94.490 177.850 ;
        RECT 94.660 177.295 94.920 178.020 ;
        RECT 95.090 177.125 95.350 177.850 ;
        RECT 95.520 177.295 95.780 178.020 ;
        RECT 95.950 177.125 96.210 177.850 ;
        RECT 96.380 177.295 96.640 178.020 ;
        RECT 96.810 177.125 97.070 177.850 ;
        RECT 97.240 177.295 97.485 178.020 ;
        RECT 97.655 177.125 97.915 177.850 ;
        RECT 98.100 177.295 98.345 178.020 ;
        RECT 98.515 177.125 98.775 177.850 ;
        RECT 98.960 177.295 99.205 178.020 ;
        RECT 99.375 177.125 99.635 177.850 ;
        RECT 99.820 177.295 100.075 178.020 ;
        RECT 94.230 177.110 99.635 177.125 ;
        RECT 100.245 177.110 100.535 177.850 ;
        RECT 100.705 177.280 100.975 178.025 ;
        RECT 94.230 176.885 100.975 177.110 ;
        RECT 84.675 175.475 90.020 176.020 ;
        RECT 90.195 175.475 91.865 176.245 ;
        RECT 92.035 176.155 92.350 176.715 ;
        RECT 92.520 176.465 99.640 176.715 ;
        RECT 92.035 175.475 92.340 175.985 ;
        RECT 92.520 175.655 92.770 176.465 ;
        RECT 92.940 175.475 93.200 176.000 ;
        RECT 93.380 175.655 93.630 176.465 ;
        RECT 99.810 176.295 100.975 176.885 ;
        RECT 94.230 176.125 100.975 176.295 ;
        RECT 101.235 176.885 101.620 177.855 ;
        RECT 101.790 177.565 102.115 178.025 ;
        RECT 102.635 177.395 102.915 177.855 ;
        RECT 101.790 177.175 102.915 177.395 ;
        RECT 101.235 176.215 101.515 176.885 ;
        RECT 101.790 176.715 102.240 177.175 ;
        RECT 103.105 177.005 103.505 177.855 ;
        RECT 103.905 177.565 104.175 178.025 ;
        RECT 104.345 177.395 104.630 177.855 ;
        RECT 101.685 176.385 102.240 176.715 ;
        RECT 102.410 176.445 103.505 177.005 ;
        RECT 101.790 176.275 102.240 176.385 ;
        RECT 93.800 175.475 94.060 176.035 ;
        RECT 94.230 175.670 94.490 176.125 ;
        RECT 94.660 175.475 94.920 175.955 ;
        RECT 95.090 175.670 95.350 176.125 ;
        RECT 95.520 175.475 95.780 175.955 ;
        RECT 95.950 175.670 96.210 176.125 ;
        RECT 96.380 175.475 96.625 175.955 ;
        RECT 96.795 175.670 97.070 176.125 ;
        RECT 97.240 175.475 97.485 175.955 ;
        RECT 97.655 175.670 97.915 176.125 ;
        RECT 98.095 175.475 98.345 175.955 ;
        RECT 98.515 175.670 98.775 176.125 ;
        RECT 98.955 175.475 99.205 175.955 ;
        RECT 99.375 175.670 99.635 176.125 ;
        RECT 99.815 175.475 100.075 175.955 ;
        RECT 100.245 175.670 100.505 176.125 ;
        RECT 100.675 175.475 100.975 175.955 ;
        RECT 101.235 175.645 101.620 176.215 ;
        RECT 101.790 176.105 102.915 176.275 ;
        RECT 101.790 175.475 102.115 175.935 ;
        RECT 102.635 175.645 102.915 176.105 ;
        RECT 103.105 175.645 103.505 176.445 ;
        RECT 103.675 177.175 104.630 177.395 ;
        RECT 103.675 176.275 103.885 177.175 ;
        RECT 104.055 176.445 104.745 177.005 ;
        RECT 105.375 176.885 105.760 177.855 ;
        RECT 105.930 177.565 106.255 178.025 ;
        RECT 106.775 177.395 107.055 177.855 ;
        RECT 105.930 177.175 107.055 177.395 ;
        RECT 103.675 176.105 104.630 176.275 ;
        RECT 103.905 175.475 104.175 175.935 ;
        RECT 104.345 175.645 104.630 176.105 ;
        RECT 105.375 176.215 105.655 176.885 ;
        RECT 105.930 176.715 106.380 177.175 ;
        RECT 107.245 177.005 107.645 177.855 ;
        RECT 108.045 177.565 108.315 178.025 ;
        RECT 108.485 177.395 108.770 177.855 ;
        RECT 105.825 176.385 106.380 176.715 ;
        RECT 106.550 176.445 107.645 177.005 ;
        RECT 105.930 176.275 106.380 176.385 ;
        RECT 105.375 175.645 105.760 176.215 ;
        RECT 105.930 176.105 107.055 176.275 ;
        RECT 105.930 175.475 106.255 175.935 ;
        RECT 106.775 175.645 107.055 176.105 ;
        RECT 107.245 175.645 107.645 176.445 ;
        RECT 107.815 177.175 108.770 177.395 ;
        RECT 107.815 176.275 108.025 177.175 ;
        RECT 108.195 176.445 108.885 177.005 ;
        RECT 109.975 176.860 110.265 178.025 ;
        RECT 110.440 176.885 110.775 177.855 ;
        RECT 110.945 176.885 111.115 178.025 ;
        RECT 111.285 177.685 113.315 177.855 ;
        RECT 107.815 176.105 108.770 176.275 ;
        RECT 110.440 176.215 110.610 176.885 ;
        RECT 111.285 176.715 111.455 177.685 ;
        RECT 110.780 176.385 111.035 176.715 ;
        RECT 111.260 176.385 111.455 176.715 ;
        RECT 111.625 177.345 112.750 177.515 ;
        RECT 110.865 176.215 111.035 176.385 ;
        RECT 111.625 176.215 111.795 177.345 ;
        RECT 108.045 175.475 108.315 175.935 ;
        RECT 108.485 175.645 108.770 176.105 ;
        RECT 109.975 175.475 110.265 176.200 ;
        RECT 110.440 175.645 110.695 176.215 ;
        RECT 110.865 176.045 111.795 176.215 ;
        RECT 111.965 177.005 112.975 177.175 ;
        RECT 111.965 176.205 112.135 177.005 ;
        RECT 112.340 176.665 112.615 176.805 ;
        RECT 112.335 176.495 112.615 176.665 ;
        RECT 111.620 176.010 111.795 176.045 ;
        RECT 110.865 175.475 111.195 175.875 ;
        RECT 111.620 175.645 112.150 176.010 ;
        RECT 112.340 175.645 112.615 176.495 ;
        RECT 112.785 175.645 112.975 177.005 ;
        RECT 113.145 177.020 113.315 177.685 ;
        RECT 113.485 177.265 113.655 178.025 ;
        RECT 113.890 177.265 114.405 177.675 ;
        RECT 113.145 176.830 113.895 177.020 ;
        RECT 114.065 176.455 114.405 177.265 ;
        RECT 114.575 176.885 114.835 178.025 ;
        RECT 115.005 176.875 115.335 177.855 ;
        RECT 115.505 176.885 115.785 178.025 ;
        RECT 115.955 176.885 116.215 178.025 ;
        RECT 116.385 176.875 116.715 177.855 ;
        RECT 116.885 176.885 117.165 178.025 ;
        RECT 118.255 176.935 119.465 178.025 ;
        RECT 114.595 176.465 114.930 176.715 ;
        RECT 113.175 176.285 114.405 176.455 ;
        RECT 113.155 175.475 113.665 176.010 ;
        RECT 113.885 175.680 114.130 176.285 ;
        RECT 115.100 176.275 115.270 176.875 ;
        RECT 115.440 176.445 115.775 176.715 ;
        RECT 115.975 176.465 116.310 176.715 ;
        RECT 116.480 176.275 116.650 176.875 ;
        RECT 116.820 176.445 117.155 176.715 ;
        RECT 118.255 176.395 118.775 176.935 ;
        RECT 114.575 175.645 115.270 176.275 ;
        RECT 115.475 175.475 115.785 176.275 ;
        RECT 115.955 175.645 116.650 176.275 ;
        RECT 116.855 175.475 117.165 176.275 ;
        RECT 118.945 176.225 119.465 176.765 ;
        RECT 118.255 175.475 119.465 176.225 ;
        RECT 71.250 175.305 119.550 175.475 ;
        RECT 71.335 174.555 72.545 175.305 ;
        RECT 72.715 174.555 73.925 175.305 ;
        RECT 74.100 174.755 74.355 175.045 ;
        RECT 74.525 174.925 74.855 175.305 ;
        RECT 74.100 174.585 74.850 174.755 ;
        RECT 71.335 174.015 71.855 174.555 ;
        RECT 72.025 173.845 72.545 174.385 ;
        RECT 72.715 174.015 73.235 174.555 ;
        RECT 73.405 173.845 73.925 174.385 ;
        RECT 71.335 172.755 72.545 173.845 ;
        RECT 72.715 172.755 73.925 173.845 ;
        RECT 74.100 173.765 74.450 174.415 ;
        RECT 74.620 173.595 74.850 174.585 ;
        RECT 74.100 173.425 74.850 173.595 ;
        RECT 74.100 172.925 74.355 173.425 ;
        RECT 74.525 172.755 74.855 173.255 ;
        RECT 75.025 172.925 75.195 175.045 ;
        RECT 75.555 174.945 75.885 175.305 ;
        RECT 76.055 174.915 76.550 175.085 ;
        RECT 76.755 174.915 77.610 175.085 ;
        RECT 75.425 173.725 75.885 174.775 ;
        RECT 75.365 172.940 75.690 173.725 ;
        RECT 76.055 173.555 76.225 174.915 ;
        RECT 76.395 174.005 76.745 174.625 ;
        RECT 76.915 174.405 77.270 174.625 ;
        RECT 76.915 173.815 77.085 174.405 ;
        RECT 77.440 174.205 77.610 174.915 ;
        RECT 78.485 174.845 78.815 175.305 ;
        RECT 79.025 174.945 79.375 175.115 ;
        RECT 77.815 174.375 78.605 174.625 ;
        RECT 79.025 174.555 79.285 174.945 ;
        RECT 79.595 174.855 80.545 175.135 ;
        RECT 80.715 174.865 80.905 175.305 ;
        RECT 81.075 174.925 82.145 175.095 ;
        RECT 78.775 174.205 78.945 174.385 ;
        RECT 76.055 173.385 76.450 173.555 ;
        RECT 76.620 173.425 77.085 173.815 ;
        RECT 77.255 174.035 78.945 174.205 ;
        RECT 76.280 173.255 76.450 173.385 ;
        RECT 77.255 173.255 77.425 174.035 ;
        RECT 79.115 173.865 79.285 174.555 ;
        RECT 77.785 173.695 79.285 173.865 ;
        RECT 79.475 173.895 79.685 174.685 ;
        RECT 79.855 174.065 80.205 174.685 ;
        RECT 80.375 174.075 80.545 174.855 ;
        RECT 81.075 174.695 81.245 174.925 ;
        RECT 80.715 174.525 81.245 174.695 ;
        RECT 80.715 174.245 80.935 174.525 ;
        RECT 81.415 174.355 81.655 174.755 ;
        RECT 80.375 173.905 80.780 174.075 ;
        RECT 81.115 173.985 81.655 174.355 ;
        RECT 81.825 174.570 82.145 174.925 ;
        RECT 82.390 174.845 82.695 175.305 ;
        RECT 82.865 174.595 83.120 175.125 ;
        RECT 81.825 174.395 82.150 174.570 ;
        RECT 81.825 174.095 82.740 174.395 ;
        RECT 82.000 174.065 82.740 174.095 ;
        RECT 79.475 173.735 80.150 173.895 ;
        RECT 80.610 173.815 80.780 173.905 ;
        RECT 79.475 173.725 80.440 173.735 ;
        RECT 79.115 173.555 79.285 173.695 ;
        RECT 75.860 172.755 76.110 173.215 ;
        RECT 76.280 172.925 76.530 173.255 ;
        RECT 76.745 172.925 77.425 173.255 ;
        RECT 77.595 173.355 78.670 173.525 ;
        RECT 79.115 173.385 79.675 173.555 ;
        RECT 79.980 173.435 80.440 173.725 ;
        RECT 80.610 173.645 81.830 173.815 ;
        RECT 77.595 173.015 77.765 173.355 ;
        RECT 78.000 172.755 78.330 173.185 ;
        RECT 78.500 173.015 78.670 173.355 ;
        RECT 78.965 172.755 79.335 173.215 ;
        RECT 79.505 172.925 79.675 173.385 ;
        RECT 80.610 173.265 80.780 173.645 ;
        RECT 82.000 173.475 82.170 174.065 ;
        RECT 82.910 173.945 83.120 174.595 ;
        RECT 83.295 174.555 84.505 175.305 ;
        RECT 84.680 174.755 84.935 175.045 ;
        RECT 85.105 174.925 85.435 175.305 ;
        RECT 84.680 174.585 85.430 174.755 ;
        RECT 83.295 174.015 83.815 174.555 ;
        RECT 79.910 172.925 80.780 173.265 ;
        RECT 81.370 173.305 82.170 173.475 ;
        RECT 80.950 172.755 81.200 173.215 ;
        RECT 81.370 173.015 81.540 173.305 ;
        RECT 81.720 172.755 82.050 173.135 ;
        RECT 82.390 172.755 82.695 173.895 ;
        RECT 82.865 173.065 83.120 173.945 ;
        RECT 83.985 173.845 84.505 174.385 ;
        RECT 83.295 172.755 84.505 173.845 ;
        RECT 84.680 173.765 85.030 174.415 ;
        RECT 85.200 173.595 85.430 174.585 ;
        RECT 84.680 173.425 85.430 173.595 ;
        RECT 84.680 172.925 84.935 173.425 ;
        RECT 85.105 172.755 85.435 173.255 ;
        RECT 85.605 172.925 85.775 175.045 ;
        RECT 86.135 174.945 86.465 175.305 ;
        RECT 86.635 174.915 87.130 175.085 ;
        RECT 87.335 174.915 88.190 175.085 ;
        RECT 86.005 173.725 86.465 174.775 ;
        RECT 85.945 172.940 86.270 173.725 ;
        RECT 86.635 173.555 86.805 174.915 ;
        RECT 86.975 174.005 87.325 174.625 ;
        RECT 87.495 174.405 87.850 174.625 ;
        RECT 87.495 173.815 87.665 174.405 ;
        RECT 88.020 174.205 88.190 174.915 ;
        RECT 89.065 174.845 89.395 175.305 ;
        RECT 89.605 174.945 89.955 175.115 ;
        RECT 88.395 174.375 89.185 174.625 ;
        RECT 89.605 174.555 89.865 174.945 ;
        RECT 90.175 174.855 91.125 175.135 ;
        RECT 91.295 174.865 91.485 175.305 ;
        RECT 91.655 174.925 92.725 175.095 ;
        RECT 89.355 174.205 89.525 174.385 ;
        RECT 86.635 173.385 87.030 173.555 ;
        RECT 87.200 173.425 87.665 173.815 ;
        RECT 87.835 174.035 89.525 174.205 ;
        RECT 86.860 173.255 87.030 173.385 ;
        RECT 87.835 173.255 88.005 174.035 ;
        RECT 89.695 173.865 89.865 174.555 ;
        RECT 88.365 173.695 89.865 173.865 ;
        RECT 90.055 173.895 90.265 174.685 ;
        RECT 90.435 174.065 90.785 174.685 ;
        RECT 90.955 174.075 91.125 174.855 ;
        RECT 91.655 174.695 91.825 174.925 ;
        RECT 91.295 174.525 91.825 174.695 ;
        RECT 91.295 174.245 91.515 174.525 ;
        RECT 91.995 174.355 92.235 174.755 ;
        RECT 90.955 173.905 91.360 174.075 ;
        RECT 91.695 173.985 92.235 174.355 ;
        RECT 92.405 174.570 92.725 174.925 ;
        RECT 92.970 174.845 93.275 175.305 ;
        RECT 93.445 174.595 93.700 175.125 ;
        RECT 92.405 174.395 92.730 174.570 ;
        RECT 92.405 174.095 93.320 174.395 ;
        RECT 92.580 174.065 93.320 174.095 ;
        RECT 90.055 173.735 90.730 173.895 ;
        RECT 91.190 173.815 91.360 173.905 ;
        RECT 90.055 173.725 91.020 173.735 ;
        RECT 89.695 173.555 89.865 173.695 ;
        RECT 86.440 172.755 86.690 173.215 ;
        RECT 86.860 172.925 87.110 173.255 ;
        RECT 87.325 172.925 88.005 173.255 ;
        RECT 88.175 173.355 89.250 173.525 ;
        RECT 89.695 173.385 90.255 173.555 ;
        RECT 90.560 173.435 91.020 173.725 ;
        RECT 91.190 173.645 92.410 173.815 ;
        RECT 88.175 173.015 88.345 173.355 ;
        RECT 88.580 172.755 88.910 173.185 ;
        RECT 89.080 173.015 89.250 173.355 ;
        RECT 89.545 172.755 89.915 173.215 ;
        RECT 90.085 172.925 90.255 173.385 ;
        RECT 91.190 173.265 91.360 173.645 ;
        RECT 92.580 173.475 92.750 174.065 ;
        RECT 93.490 173.945 93.700 174.595 ;
        RECT 90.490 172.925 91.360 173.265 ;
        RECT 91.950 173.305 92.750 173.475 ;
        RECT 91.530 172.755 91.780 173.215 ;
        RECT 91.950 173.015 92.120 173.305 ;
        RECT 92.300 172.755 92.630 173.135 ;
        RECT 92.970 172.755 93.275 173.895 ;
        RECT 93.445 173.065 93.700 173.945 ;
        RECT 94.335 174.360 94.675 175.135 ;
        RECT 94.845 174.845 95.015 175.305 ;
        RECT 95.255 174.870 95.615 175.135 ;
        RECT 95.255 174.865 95.610 174.870 ;
        RECT 95.255 174.855 95.605 174.865 ;
        RECT 95.255 174.850 95.600 174.855 ;
        RECT 95.255 174.840 95.595 174.850 ;
        RECT 96.245 174.845 96.415 175.305 ;
        RECT 95.255 174.835 95.590 174.840 ;
        RECT 95.255 174.825 95.580 174.835 ;
        RECT 95.255 174.815 95.570 174.825 ;
        RECT 95.255 174.675 95.555 174.815 ;
        RECT 94.845 174.485 95.555 174.675 ;
        RECT 95.745 174.675 96.075 174.755 ;
        RECT 96.585 174.675 96.925 175.135 ;
        RECT 95.745 174.485 96.925 174.675 ;
        RECT 97.095 174.580 97.385 175.305 ;
        RECT 97.645 174.755 97.815 175.045 ;
        RECT 97.985 174.925 98.315 175.305 ;
        RECT 97.645 174.585 98.310 174.755 ;
        RECT 94.335 172.925 94.615 174.360 ;
        RECT 94.845 173.915 95.130 174.485 ;
        RECT 95.315 174.085 95.785 174.315 ;
        RECT 95.955 174.295 96.285 174.315 ;
        RECT 95.955 174.115 96.405 174.295 ;
        RECT 96.595 174.115 96.925 174.315 ;
        RECT 94.845 173.700 95.995 173.915 ;
        RECT 94.785 172.755 95.495 173.530 ;
        RECT 95.665 172.925 95.995 173.700 ;
        RECT 96.190 173.000 96.405 174.115 ;
        RECT 96.695 173.775 96.925 174.115 ;
        RECT 96.585 172.755 96.915 173.475 ;
        RECT 97.095 172.755 97.385 173.920 ;
        RECT 97.560 173.765 97.910 174.415 ;
        RECT 98.080 173.595 98.310 174.585 ;
        RECT 97.645 173.425 98.310 173.595 ;
        RECT 97.645 172.925 97.815 173.425 ;
        RECT 97.985 172.755 98.315 173.255 ;
        RECT 98.485 172.925 98.670 175.045 ;
        RECT 98.925 174.845 99.175 175.305 ;
        RECT 99.345 174.855 99.680 175.025 ;
        RECT 99.875 174.855 100.550 175.025 ;
        RECT 99.345 174.715 99.515 174.855 ;
        RECT 98.840 173.725 99.120 174.675 ;
        RECT 99.290 174.585 99.515 174.715 ;
        RECT 99.290 173.480 99.460 174.585 ;
        RECT 99.685 174.435 100.210 174.655 ;
        RECT 99.630 173.670 99.870 174.265 ;
        RECT 100.040 173.735 100.210 174.435 ;
        RECT 100.380 174.075 100.550 174.855 ;
        RECT 100.870 174.805 101.240 175.305 ;
        RECT 101.420 174.855 101.825 175.025 ;
        RECT 101.995 174.855 102.780 175.025 ;
        RECT 101.420 174.625 101.590 174.855 ;
        RECT 100.760 174.325 101.590 174.625 ;
        RECT 101.975 174.355 102.440 174.685 ;
        RECT 100.760 174.295 100.960 174.325 ;
        RECT 101.080 174.075 101.250 174.145 ;
        RECT 100.380 173.905 101.250 174.075 ;
        RECT 100.740 173.815 101.250 173.905 ;
        RECT 99.290 173.350 99.595 173.480 ;
        RECT 100.040 173.370 100.570 173.735 ;
        RECT 98.910 172.755 99.175 173.215 ;
        RECT 99.345 172.925 99.595 173.350 ;
        RECT 100.740 173.200 100.910 173.815 ;
        RECT 99.805 173.030 100.910 173.200 ;
        RECT 101.080 172.755 101.250 173.555 ;
        RECT 101.420 173.255 101.590 174.325 ;
        RECT 101.760 173.425 101.950 174.145 ;
        RECT 102.120 173.395 102.440 174.355 ;
        RECT 102.610 174.395 102.780 174.855 ;
        RECT 103.055 174.775 103.265 175.305 ;
        RECT 103.525 174.565 103.855 175.090 ;
        RECT 104.025 174.695 104.195 175.305 ;
        RECT 104.365 174.650 104.695 175.085 ;
        RECT 104.365 174.565 104.745 174.650 ;
        RECT 103.655 174.395 103.855 174.565 ;
        RECT 104.520 174.525 104.745 174.565 ;
        RECT 102.610 174.065 103.485 174.395 ;
        RECT 103.655 174.065 104.405 174.395 ;
        RECT 101.420 172.925 101.670 173.255 ;
        RECT 102.610 173.225 102.780 174.065 ;
        RECT 103.655 173.860 103.845 174.065 ;
        RECT 104.575 173.945 104.745 174.525 ;
        RECT 105.650 174.495 105.895 175.100 ;
        RECT 106.115 174.770 106.625 175.305 ;
        RECT 104.530 173.895 104.745 173.945 ;
        RECT 102.950 173.485 103.845 173.860 ;
        RECT 104.355 173.815 104.745 173.895 ;
        RECT 105.375 174.325 106.605 174.495 ;
        RECT 101.895 173.055 102.780 173.225 ;
        RECT 102.960 172.755 103.275 173.255 ;
        RECT 103.505 172.925 103.845 173.485 ;
        RECT 104.015 172.755 104.185 173.765 ;
        RECT 104.355 172.970 104.685 173.815 ;
        RECT 105.375 173.515 105.715 174.325 ;
        RECT 105.885 173.760 106.635 173.950 ;
        RECT 105.375 173.105 105.890 173.515 ;
        RECT 106.125 172.755 106.295 173.515 ;
        RECT 106.465 173.095 106.635 173.760 ;
        RECT 106.805 173.775 106.995 175.135 ;
        RECT 107.165 174.965 107.440 175.135 ;
        RECT 107.165 174.795 107.445 174.965 ;
        RECT 107.165 173.975 107.440 174.795 ;
        RECT 107.630 174.770 108.160 175.135 ;
        RECT 108.585 174.905 108.915 175.305 ;
        RECT 107.985 174.735 108.160 174.770 ;
        RECT 107.645 173.775 107.815 174.575 ;
        RECT 106.805 173.605 107.815 173.775 ;
        RECT 107.985 174.565 108.915 174.735 ;
        RECT 109.085 174.565 109.340 175.135 ;
        RECT 107.985 173.435 108.155 174.565 ;
        RECT 108.745 174.395 108.915 174.565 ;
        RECT 107.030 173.265 108.155 173.435 ;
        RECT 108.325 174.065 108.520 174.395 ;
        RECT 108.745 174.065 109.000 174.395 ;
        RECT 108.325 173.095 108.495 174.065 ;
        RECT 109.170 173.895 109.340 174.565 ;
        RECT 109.525 174.495 109.795 175.305 ;
        RECT 109.965 174.495 110.295 175.135 ;
        RECT 110.465 174.495 110.705 175.305 ;
        RECT 111.630 174.495 111.875 175.100 ;
        RECT 112.095 174.770 112.605 175.305 ;
        RECT 109.515 174.065 109.865 174.315 ;
        RECT 110.035 173.895 110.205 174.495 ;
        RECT 111.355 174.325 112.585 174.495 ;
        RECT 110.375 174.065 110.725 174.315 ;
        RECT 106.465 172.925 108.495 173.095 ;
        RECT 108.665 172.755 108.835 173.895 ;
        RECT 109.005 172.925 109.340 173.895 ;
        RECT 109.525 172.755 109.855 173.895 ;
        RECT 110.035 173.725 110.715 173.895 ;
        RECT 110.385 172.940 110.715 173.725 ;
        RECT 111.355 173.515 111.695 174.325 ;
        RECT 111.865 173.760 112.615 173.950 ;
        RECT 111.355 173.105 111.870 173.515 ;
        RECT 112.105 172.755 112.275 173.515 ;
        RECT 112.445 173.095 112.615 173.760 ;
        RECT 112.785 173.775 112.975 175.135 ;
        RECT 113.145 174.965 113.420 175.135 ;
        RECT 113.145 174.795 113.425 174.965 ;
        RECT 113.145 173.975 113.420 174.795 ;
        RECT 113.610 174.770 114.140 175.135 ;
        RECT 114.565 174.905 114.895 175.305 ;
        RECT 113.965 174.735 114.140 174.770 ;
        RECT 113.625 173.775 113.795 174.575 ;
        RECT 112.785 173.605 113.795 173.775 ;
        RECT 113.965 174.565 114.895 174.735 ;
        RECT 115.065 174.565 115.320 175.135 ;
        RECT 113.965 173.435 114.135 174.565 ;
        RECT 114.725 174.395 114.895 174.565 ;
        RECT 113.010 173.265 114.135 173.435 ;
        RECT 114.305 174.065 114.500 174.395 ;
        RECT 114.725 174.065 114.980 174.395 ;
        RECT 114.305 173.095 114.475 174.065 ;
        RECT 115.150 173.895 115.320 174.565 ;
        RECT 112.445 172.925 114.475 173.095 ;
        RECT 114.645 172.755 114.815 173.895 ;
        RECT 114.985 172.925 115.320 173.895 ;
        RECT 115.530 174.565 116.145 175.135 ;
        RECT 116.315 174.795 116.530 175.305 ;
        RECT 116.760 174.795 117.040 175.125 ;
        RECT 117.220 174.795 117.460 175.305 ;
        RECT 115.530 173.545 115.845 174.565 ;
        RECT 116.015 173.895 116.185 174.395 ;
        RECT 116.435 174.065 116.700 174.625 ;
        RECT 116.870 173.895 117.040 174.795 ;
        RECT 117.210 174.065 117.565 174.625 ;
        RECT 118.255 174.555 119.465 175.305 ;
        RECT 116.015 173.725 117.440 173.895 ;
        RECT 115.530 172.925 116.065 173.545 ;
        RECT 116.235 172.755 116.565 173.555 ;
        RECT 117.050 173.550 117.440 173.725 ;
        RECT 118.255 173.845 118.775 174.385 ;
        RECT 118.945 174.015 119.465 174.555 ;
        RECT 118.255 172.755 119.465 173.845 ;
        RECT 71.250 172.585 119.550 172.755 ;
        RECT 71.335 171.495 72.545 172.585 ;
        RECT 72.715 171.495 74.385 172.585 ;
        RECT 75.035 172.075 75.335 172.585 ;
        RECT 75.505 172.075 75.885 172.245 ;
        RECT 76.465 172.075 77.095 172.585 ;
        RECT 75.505 171.905 75.675 172.075 ;
        RECT 77.265 171.905 77.595 172.415 ;
        RECT 77.765 172.075 78.065 172.585 ;
        RECT 78.235 172.150 83.580 172.585 ;
        RECT 71.335 170.785 71.855 171.325 ;
        RECT 72.025 170.955 72.545 171.495 ;
        RECT 72.715 170.805 73.465 171.325 ;
        RECT 73.635 170.975 74.385 171.495 ;
        RECT 75.015 171.705 75.675 171.905 ;
        RECT 75.845 171.735 78.065 171.905 ;
        RECT 71.335 170.035 72.545 170.785 ;
        RECT 72.715 170.035 74.385 170.805 ;
        RECT 75.015 170.775 75.185 171.705 ;
        RECT 75.845 171.535 76.015 171.735 ;
        RECT 75.355 171.365 76.015 171.535 ;
        RECT 76.185 171.395 77.725 171.565 ;
        RECT 75.355 170.945 75.525 171.365 ;
        RECT 76.185 171.195 76.355 171.395 ;
        RECT 75.755 171.025 76.355 171.195 ;
        RECT 76.525 171.025 77.220 171.225 ;
        RECT 77.480 170.945 77.725 171.395 ;
        RECT 75.845 170.775 76.755 170.855 ;
        RECT 75.015 170.295 75.335 170.775 ;
        RECT 75.505 170.685 76.755 170.775 ;
        RECT 75.505 170.605 76.015 170.685 ;
        RECT 75.505 170.205 75.735 170.605 ;
        RECT 75.905 170.035 76.255 170.425 ;
        RECT 76.425 170.205 76.755 170.685 ;
        RECT 76.925 170.035 77.095 170.855 ;
        RECT 77.895 170.775 78.065 171.735 ;
        RECT 77.600 170.230 78.065 170.775 ;
        RECT 79.820 170.580 80.160 171.410 ;
        RECT 81.640 170.900 81.990 172.150 ;
        RECT 84.215 171.420 84.505 172.585 ;
        RECT 84.755 171.655 84.935 172.415 ;
        RECT 85.115 171.825 85.445 172.585 ;
        RECT 84.755 171.485 85.430 171.655 ;
        RECT 85.615 171.510 85.885 172.415 ;
        RECT 85.260 171.340 85.430 171.485 ;
        RECT 84.695 170.935 85.035 171.305 ;
        RECT 85.260 171.010 85.535 171.340 ;
        RECT 78.235 170.035 83.580 170.580 ;
        RECT 84.215 170.035 84.505 170.760 ;
        RECT 85.260 170.755 85.430 171.010 ;
        RECT 84.765 170.585 85.430 170.755 ;
        RECT 85.705 170.710 85.885 171.510 ;
        RECT 86.055 171.495 87.725 172.585 ;
        RECT 84.765 170.205 84.935 170.585 ;
        RECT 85.115 170.035 85.445 170.415 ;
        RECT 85.625 170.205 85.885 170.710 ;
        RECT 86.055 170.805 86.805 171.325 ;
        RECT 86.975 170.975 87.725 171.495 ;
        RECT 87.895 171.445 88.155 172.415 ;
        RECT 88.325 172.160 88.710 172.585 ;
        RECT 88.880 171.990 89.135 172.415 ;
        RECT 88.325 171.795 89.135 171.990 ;
        RECT 86.055 170.035 87.725 170.805 ;
        RECT 87.895 170.775 88.080 171.445 ;
        RECT 88.325 171.275 88.675 171.795 ;
        RECT 89.325 171.625 89.570 172.415 ;
        RECT 89.740 172.160 90.125 172.585 ;
        RECT 90.295 171.990 90.570 172.415 ;
        RECT 88.250 170.945 88.675 171.275 ;
        RECT 88.845 171.445 89.570 171.625 ;
        RECT 89.740 171.795 90.570 171.990 ;
        RECT 88.845 170.945 89.495 171.445 ;
        RECT 89.740 171.275 90.090 171.795 ;
        RECT 90.740 171.625 91.165 172.415 ;
        RECT 91.335 172.160 91.720 172.585 ;
        RECT 91.890 171.990 92.325 172.415 ;
        RECT 89.665 170.945 90.090 171.275 ;
        RECT 90.260 171.445 91.165 171.625 ;
        RECT 91.335 171.820 92.325 171.990 ;
        RECT 90.260 170.945 91.090 171.445 ;
        RECT 91.335 171.275 91.670 171.820 ;
        RECT 92.505 171.775 92.800 172.585 ;
        RECT 91.260 170.945 91.670 171.275 ;
        RECT 91.840 170.945 92.325 171.650 ;
        RECT 92.980 171.275 93.225 172.415 ;
        RECT 93.400 171.775 93.660 172.585 ;
        RECT 94.260 172.580 100.535 172.585 ;
        RECT 93.840 171.275 94.090 172.410 ;
        RECT 94.260 171.785 94.520 172.580 ;
        RECT 94.690 171.685 94.950 172.410 ;
        RECT 95.120 171.855 95.380 172.580 ;
        RECT 95.550 171.685 95.810 172.410 ;
        RECT 95.980 171.855 96.240 172.580 ;
        RECT 96.410 171.685 96.670 172.410 ;
        RECT 96.840 171.855 97.100 172.580 ;
        RECT 97.270 171.685 97.530 172.410 ;
        RECT 97.700 171.855 97.945 172.580 ;
        RECT 98.115 171.685 98.375 172.410 ;
        RECT 98.560 171.855 98.805 172.580 ;
        RECT 98.975 171.685 99.235 172.410 ;
        RECT 99.420 171.855 99.665 172.580 ;
        RECT 99.835 171.685 100.095 172.410 ;
        RECT 100.280 171.855 100.535 172.580 ;
        RECT 94.690 171.670 100.095 171.685 ;
        RECT 100.705 171.670 100.995 172.410 ;
        RECT 101.165 171.840 101.435 172.585 ;
        RECT 102.705 171.915 102.875 172.415 ;
        RECT 103.045 172.085 103.375 172.585 ;
        RECT 102.705 171.745 103.370 171.915 ;
        RECT 94.690 171.445 101.435 171.670 ;
        RECT 88.325 170.775 88.675 170.945 ;
        RECT 89.325 170.775 89.495 170.945 ;
        RECT 89.740 170.775 90.090 170.945 ;
        RECT 90.740 170.775 91.090 170.945 ;
        RECT 91.335 170.775 91.670 170.945 ;
        RECT 87.895 170.205 88.155 170.775 ;
        RECT 88.325 170.605 89.135 170.775 ;
        RECT 88.325 170.035 88.710 170.435 ;
        RECT 88.880 170.205 89.135 170.605 ;
        RECT 89.325 170.205 89.570 170.775 ;
        RECT 89.740 170.605 90.550 170.775 ;
        RECT 89.740 170.035 90.125 170.435 ;
        RECT 90.295 170.205 90.550 170.605 ;
        RECT 90.740 170.205 91.165 170.775 ;
        RECT 91.335 170.605 92.325 170.775 ;
        RECT 92.495 170.715 92.810 171.275 ;
        RECT 92.980 171.025 100.100 171.275 ;
        RECT 91.335 170.035 91.720 170.435 ;
        RECT 91.890 170.205 92.325 170.605 ;
        RECT 92.495 170.035 92.800 170.545 ;
        RECT 92.980 170.215 93.230 171.025 ;
        RECT 93.400 170.035 93.660 170.560 ;
        RECT 93.840 170.215 94.090 171.025 ;
        RECT 100.270 170.855 101.435 171.445 ;
        RECT 102.620 170.925 102.970 171.575 ;
        RECT 94.690 170.685 101.435 170.855 ;
        RECT 103.140 170.755 103.370 171.745 ;
        RECT 94.260 170.035 94.520 170.595 ;
        RECT 94.690 170.230 94.950 170.685 ;
        RECT 95.120 170.035 95.380 170.515 ;
        RECT 95.550 170.230 95.810 170.685 ;
        RECT 95.980 170.035 96.240 170.515 ;
        RECT 96.410 170.230 96.670 170.685 ;
        RECT 96.840 170.035 97.085 170.515 ;
        RECT 97.255 170.230 97.530 170.685 ;
        RECT 97.700 170.035 97.945 170.515 ;
        RECT 98.115 170.230 98.375 170.685 ;
        RECT 98.555 170.035 98.805 170.515 ;
        RECT 98.975 170.230 99.235 170.685 ;
        RECT 99.415 170.035 99.665 170.515 ;
        RECT 99.835 170.230 100.095 170.685 ;
        RECT 100.275 170.035 100.535 170.515 ;
        RECT 100.705 170.230 100.965 170.685 ;
        RECT 102.705 170.585 103.370 170.755 ;
        RECT 101.135 170.035 101.435 170.515 ;
        RECT 102.705 170.295 102.875 170.585 ;
        RECT 103.045 170.035 103.375 170.415 ;
        RECT 103.545 170.295 103.730 172.415 ;
        RECT 103.970 172.125 104.235 172.585 ;
        RECT 104.405 171.990 104.655 172.415 ;
        RECT 104.865 172.140 105.970 172.310 ;
        RECT 104.350 171.860 104.655 171.990 ;
        RECT 103.900 170.665 104.180 171.615 ;
        RECT 104.350 170.755 104.520 171.860 ;
        RECT 104.690 171.075 104.930 171.670 ;
        RECT 105.100 171.605 105.630 171.970 ;
        RECT 105.100 170.905 105.270 171.605 ;
        RECT 105.800 171.525 105.970 172.140 ;
        RECT 106.140 171.785 106.310 172.585 ;
        RECT 106.480 172.085 106.730 172.415 ;
        RECT 106.955 172.115 107.840 172.285 ;
        RECT 105.800 171.435 106.310 171.525 ;
        RECT 104.350 170.625 104.575 170.755 ;
        RECT 104.745 170.685 105.270 170.905 ;
        RECT 105.440 171.265 106.310 171.435 ;
        RECT 103.985 170.035 104.235 170.495 ;
        RECT 104.405 170.485 104.575 170.625 ;
        RECT 105.440 170.485 105.610 171.265 ;
        RECT 106.140 171.195 106.310 171.265 ;
        RECT 105.820 171.015 106.020 171.045 ;
        RECT 106.480 171.015 106.650 172.085 ;
        RECT 106.820 171.195 107.010 171.915 ;
        RECT 105.820 170.715 106.650 171.015 ;
        RECT 107.180 170.985 107.500 171.945 ;
        RECT 104.405 170.315 104.740 170.485 ;
        RECT 104.935 170.315 105.610 170.485 ;
        RECT 105.930 170.035 106.300 170.535 ;
        RECT 106.480 170.485 106.650 170.715 ;
        RECT 107.035 170.655 107.500 170.985 ;
        RECT 107.670 171.275 107.840 172.115 ;
        RECT 108.020 172.085 108.335 172.585 ;
        RECT 108.565 171.855 108.905 172.415 ;
        RECT 108.010 171.480 108.905 171.855 ;
        RECT 109.075 171.575 109.245 172.585 ;
        RECT 108.715 171.275 108.905 171.480 ;
        RECT 109.415 171.525 109.745 172.370 ;
        RECT 109.415 171.445 109.805 171.525 ;
        RECT 109.590 171.395 109.805 171.445 ;
        RECT 109.975 171.420 110.265 172.585 ;
        RECT 110.435 171.445 110.820 172.415 ;
        RECT 110.990 172.125 111.315 172.585 ;
        RECT 111.835 171.955 112.115 172.415 ;
        RECT 110.990 171.735 112.115 171.955 ;
        RECT 107.670 170.945 108.545 171.275 ;
        RECT 108.715 170.945 109.465 171.275 ;
        RECT 107.670 170.485 107.840 170.945 ;
        RECT 108.715 170.775 108.915 170.945 ;
        RECT 109.635 170.815 109.805 171.395 ;
        RECT 109.580 170.775 109.805 170.815 ;
        RECT 106.480 170.315 106.885 170.485 ;
        RECT 107.055 170.315 107.840 170.485 ;
        RECT 108.115 170.035 108.325 170.565 ;
        RECT 108.585 170.250 108.915 170.775 ;
        RECT 109.425 170.690 109.805 170.775 ;
        RECT 110.435 170.775 110.715 171.445 ;
        RECT 110.990 171.275 111.440 171.735 ;
        RECT 112.305 171.565 112.705 172.415 ;
        RECT 113.105 172.125 113.375 172.585 ;
        RECT 113.545 171.955 113.830 172.415 ;
        RECT 110.885 170.945 111.440 171.275 ;
        RECT 111.610 171.005 112.705 171.565 ;
        RECT 110.990 170.835 111.440 170.945 ;
        RECT 109.085 170.035 109.255 170.645 ;
        RECT 109.425 170.255 109.755 170.690 ;
        RECT 109.975 170.035 110.265 170.760 ;
        RECT 110.435 170.205 110.820 170.775 ;
        RECT 110.990 170.665 112.115 170.835 ;
        RECT 110.990 170.035 111.315 170.495 ;
        RECT 111.835 170.205 112.115 170.665 ;
        RECT 112.305 170.205 112.705 171.005 ;
        RECT 112.875 171.735 113.830 171.955 ;
        RECT 112.875 170.835 113.085 171.735 ;
        RECT 113.255 171.005 113.945 171.565 ;
        RECT 114.115 171.445 114.500 172.415 ;
        RECT 114.670 172.125 114.995 172.585 ;
        RECT 115.515 171.955 115.795 172.415 ;
        RECT 114.670 171.735 115.795 171.955 ;
        RECT 112.875 170.665 113.830 170.835 ;
        RECT 113.105 170.035 113.375 170.495 ;
        RECT 113.545 170.205 113.830 170.665 ;
        RECT 114.115 170.775 114.395 171.445 ;
        RECT 114.670 171.275 115.120 171.735 ;
        RECT 115.985 171.565 116.385 172.415 ;
        RECT 116.785 172.125 117.055 172.585 ;
        RECT 117.225 171.955 117.510 172.415 ;
        RECT 114.565 170.945 115.120 171.275 ;
        RECT 115.290 171.005 116.385 171.565 ;
        RECT 114.670 170.835 115.120 170.945 ;
        RECT 114.115 170.205 114.500 170.775 ;
        RECT 114.670 170.665 115.795 170.835 ;
        RECT 114.670 170.035 114.995 170.495 ;
        RECT 115.515 170.205 115.795 170.665 ;
        RECT 115.985 170.205 116.385 171.005 ;
        RECT 116.555 171.735 117.510 171.955 ;
        RECT 116.555 170.835 116.765 171.735 ;
        RECT 116.935 171.005 117.625 171.565 ;
        RECT 118.255 171.495 119.465 172.585 ;
        RECT 118.255 170.955 118.775 171.495 ;
        RECT 116.555 170.665 117.510 170.835 ;
        RECT 118.945 170.785 119.465 171.325 ;
        RECT 116.785 170.035 117.055 170.495 ;
        RECT 117.225 170.205 117.510 170.665 ;
        RECT 118.255 170.035 119.465 170.785 ;
        RECT 71.250 169.865 119.550 170.035 ;
        RECT 71.335 169.115 72.545 169.865 ;
        RECT 72.715 169.320 78.060 169.865 ;
        RECT 78.235 169.320 83.580 169.865 ;
        RECT 84.725 169.475 85.055 169.865 ;
        RECT 71.335 168.575 71.855 169.115 ;
        RECT 72.025 168.405 72.545 168.945 ;
        RECT 74.300 168.490 74.640 169.320 ;
        RECT 71.335 167.315 72.545 168.405 ;
        RECT 76.120 167.750 76.470 169.000 ;
        RECT 79.820 168.490 80.160 169.320 ;
        RECT 85.225 169.295 85.395 169.615 ;
        RECT 85.565 169.475 85.895 169.865 ;
        RECT 86.310 169.465 87.265 169.635 ;
        RECT 84.675 169.125 86.925 169.295 ;
        RECT 81.640 167.750 81.990 169.000 ;
        RECT 84.675 168.165 84.845 169.125 ;
        RECT 85.015 168.505 85.260 168.955 ;
        RECT 85.430 168.675 85.980 168.875 ;
        RECT 86.150 168.705 86.525 168.875 ;
        RECT 86.150 168.505 86.320 168.705 ;
        RECT 86.695 168.625 86.925 169.125 ;
        RECT 85.015 168.335 86.320 168.505 ;
        RECT 87.095 168.585 87.265 169.465 ;
        RECT 87.435 169.030 87.725 169.865 ;
        RECT 87.945 169.475 88.275 169.865 ;
        RECT 88.445 169.295 88.615 169.615 ;
        RECT 88.785 169.475 89.115 169.865 ;
        RECT 89.530 169.465 90.485 169.635 ;
        RECT 87.895 169.125 90.145 169.295 ;
        RECT 87.095 168.415 87.725 168.585 ;
        RECT 72.715 167.315 78.060 167.750 ;
        RECT 78.235 167.315 83.580 167.750 ;
        RECT 84.675 167.485 85.055 168.165 ;
        RECT 85.645 167.315 85.815 168.165 ;
        RECT 85.985 167.995 87.225 168.165 ;
        RECT 85.985 167.485 86.315 167.995 ;
        RECT 86.485 167.315 86.655 167.825 ;
        RECT 86.825 167.485 87.225 167.995 ;
        RECT 87.405 167.485 87.725 168.415 ;
        RECT 87.895 168.165 88.065 169.125 ;
        RECT 88.235 168.505 88.480 168.955 ;
        RECT 88.650 168.675 89.200 168.875 ;
        RECT 89.370 168.705 89.745 168.875 ;
        RECT 89.370 168.505 89.540 168.705 ;
        RECT 89.915 168.625 90.145 169.125 ;
        RECT 88.235 168.335 89.540 168.505 ;
        RECT 90.315 168.585 90.485 169.465 ;
        RECT 90.655 169.030 90.945 169.865 ;
        RECT 91.230 169.235 91.515 169.695 ;
        RECT 91.685 169.405 91.955 169.865 ;
        RECT 91.230 169.065 92.185 169.235 ;
        RECT 90.315 168.415 90.945 168.585 ;
        RECT 87.895 167.485 88.275 168.165 ;
        RECT 88.865 167.315 89.035 168.165 ;
        RECT 89.205 167.995 90.445 168.165 ;
        RECT 89.205 167.485 89.535 167.995 ;
        RECT 89.705 167.315 89.875 167.825 ;
        RECT 90.045 167.485 90.445 167.995 ;
        RECT 90.625 167.485 90.945 168.415 ;
        RECT 91.115 168.335 91.805 168.895 ;
        RECT 91.975 168.165 92.185 169.065 ;
        RECT 91.230 167.945 92.185 168.165 ;
        RECT 92.355 168.895 92.755 169.695 ;
        RECT 92.945 169.235 93.225 169.695 ;
        RECT 93.745 169.405 94.070 169.865 ;
        RECT 92.945 169.065 94.070 169.235 ;
        RECT 94.240 169.125 94.625 169.695 ;
        RECT 93.620 168.955 94.070 169.065 ;
        RECT 92.355 168.335 93.450 168.895 ;
        RECT 93.620 168.625 94.175 168.955 ;
        RECT 91.230 167.485 91.515 167.945 ;
        RECT 91.685 167.315 91.955 167.775 ;
        RECT 92.355 167.485 92.755 168.335 ;
        RECT 93.620 168.165 94.070 168.625 ;
        RECT 94.345 168.455 94.625 169.125 ;
        RECT 94.795 169.095 96.465 169.865 ;
        RECT 97.095 169.140 97.385 169.865 ;
        RECT 97.645 169.315 97.815 169.695 ;
        RECT 98.030 169.485 98.360 169.865 ;
        RECT 97.645 169.145 98.360 169.315 ;
        RECT 94.795 168.575 95.545 169.095 ;
        RECT 92.945 167.945 94.070 168.165 ;
        RECT 92.945 167.485 93.225 167.945 ;
        RECT 93.745 167.315 94.070 167.775 ;
        RECT 94.240 167.485 94.625 168.455 ;
        RECT 95.715 168.405 96.465 168.925 ;
        RECT 97.555 168.595 97.910 168.965 ;
        RECT 98.190 168.955 98.360 169.145 ;
        RECT 98.530 169.120 98.785 169.695 ;
        RECT 98.190 168.625 98.445 168.955 ;
        RECT 94.795 167.315 96.465 168.405 ;
        RECT 97.095 167.315 97.385 168.480 ;
        RECT 98.190 168.415 98.360 168.625 ;
        RECT 97.645 168.245 98.360 168.415 ;
        RECT 98.615 168.390 98.785 169.120 ;
        RECT 98.960 169.025 99.220 169.865 ;
        RECT 99.395 169.095 102.905 169.865 ;
        RECT 103.075 169.115 104.285 169.865 ;
        RECT 104.455 169.190 104.715 169.695 ;
        RECT 104.895 169.485 105.225 169.865 ;
        RECT 105.405 169.315 105.575 169.695 ;
        RECT 99.395 168.575 101.045 169.095 ;
        RECT 97.645 167.485 97.815 168.245 ;
        RECT 98.030 167.315 98.360 168.075 ;
        RECT 98.530 167.485 98.785 168.390 ;
        RECT 98.960 167.315 99.220 168.465 ;
        RECT 101.215 168.405 102.905 168.925 ;
        RECT 103.075 168.575 103.595 169.115 ;
        RECT 103.765 168.405 104.285 168.945 ;
        RECT 99.395 167.315 102.905 168.405 ;
        RECT 103.075 167.315 104.285 168.405 ;
        RECT 104.455 168.390 104.625 169.190 ;
        RECT 104.910 169.145 105.575 169.315 ;
        RECT 104.910 168.890 105.080 169.145 ;
        RECT 105.835 169.095 107.505 169.865 ;
        RECT 107.675 169.125 108.140 169.670 ;
        RECT 104.795 168.560 105.080 168.890 ;
        RECT 105.315 168.595 105.645 168.965 ;
        RECT 105.835 168.575 106.585 169.095 ;
        RECT 104.910 168.415 105.080 168.560 ;
        RECT 104.455 167.485 104.725 168.390 ;
        RECT 104.910 168.245 105.575 168.415 ;
        RECT 106.755 168.405 107.505 168.925 ;
        RECT 104.895 167.315 105.225 168.075 ;
        RECT 105.405 167.485 105.575 168.245 ;
        RECT 105.835 167.315 107.505 168.405 ;
        RECT 107.675 168.165 107.845 169.125 ;
        RECT 108.645 169.045 108.815 169.865 ;
        RECT 108.985 169.215 109.315 169.695 ;
        RECT 109.485 169.475 109.835 169.865 ;
        RECT 110.005 169.295 110.235 169.695 ;
        RECT 109.725 169.215 110.235 169.295 ;
        RECT 108.985 169.125 110.235 169.215 ;
        RECT 110.405 169.125 110.725 169.605 ;
        RECT 110.985 169.315 111.155 169.605 ;
        RECT 111.325 169.485 111.655 169.865 ;
        RECT 110.985 169.145 111.650 169.315 ;
        RECT 108.985 169.045 109.895 169.125 ;
        RECT 108.015 168.505 108.260 168.955 ;
        RECT 108.520 168.675 109.215 168.875 ;
        RECT 109.385 168.705 109.985 168.875 ;
        RECT 109.385 168.505 109.555 168.705 ;
        RECT 110.215 168.535 110.385 168.955 ;
        RECT 108.015 168.335 109.555 168.505 ;
        RECT 109.725 168.365 110.385 168.535 ;
        RECT 109.725 168.165 109.895 168.365 ;
        RECT 110.555 168.195 110.725 169.125 ;
        RECT 110.900 168.325 111.250 168.975 ;
        RECT 107.675 167.995 109.895 168.165 ;
        RECT 110.065 167.995 110.725 168.195 ;
        RECT 111.420 168.155 111.650 169.145 ;
        RECT 107.675 167.315 107.975 167.825 ;
        RECT 108.145 167.485 108.475 167.995 ;
        RECT 110.065 167.825 110.235 167.995 ;
        RECT 110.985 167.985 111.650 168.155 ;
        RECT 108.645 167.315 109.275 167.825 ;
        RECT 109.855 167.655 110.235 167.825 ;
        RECT 110.405 167.315 110.705 167.825 ;
        RECT 110.985 167.485 111.155 167.985 ;
        RECT 111.325 167.315 111.655 167.815 ;
        RECT 111.825 167.485 112.010 169.605 ;
        RECT 112.265 169.405 112.515 169.865 ;
        RECT 112.685 169.415 113.020 169.585 ;
        RECT 113.215 169.415 113.890 169.585 ;
        RECT 112.685 169.275 112.855 169.415 ;
        RECT 112.180 168.285 112.460 169.235 ;
        RECT 112.630 169.145 112.855 169.275 ;
        RECT 112.630 168.040 112.800 169.145 ;
        RECT 113.025 168.995 113.550 169.215 ;
        RECT 112.970 168.230 113.210 168.825 ;
        RECT 113.380 168.295 113.550 168.995 ;
        RECT 113.720 168.635 113.890 169.415 ;
        RECT 114.210 169.365 114.580 169.865 ;
        RECT 114.760 169.415 115.165 169.585 ;
        RECT 115.335 169.415 116.120 169.585 ;
        RECT 114.760 169.185 114.930 169.415 ;
        RECT 114.100 168.885 114.930 169.185 ;
        RECT 115.315 168.915 115.780 169.245 ;
        RECT 114.100 168.855 114.300 168.885 ;
        RECT 114.420 168.635 114.590 168.705 ;
        RECT 113.720 168.465 114.590 168.635 ;
        RECT 114.080 168.375 114.590 168.465 ;
        RECT 112.630 167.910 112.935 168.040 ;
        RECT 113.380 167.930 113.910 168.295 ;
        RECT 112.250 167.315 112.515 167.775 ;
        RECT 112.685 167.485 112.935 167.910 ;
        RECT 114.080 167.760 114.250 168.375 ;
        RECT 113.145 167.590 114.250 167.760 ;
        RECT 114.420 167.315 114.590 168.115 ;
        RECT 114.760 167.815 114.930 168.885 ;
        RECT 115.100 167.985 115.290 168.705 ;
        RECT 115.460 167.955 115.780 168.915 ;
        RECT 115.950 168.955 116.120 169.415 ;
        RECT 116.395 169.335 116.605 169.865 ;
        RECT 116.865 169.125 117.195 169.650 ;
        RECT 117.365 169.255 117.535 169.865 ;
        RECT 117.705 169.210 118.035 169.645 ;
        RECT 117.705 169.125 118.085 169.210 ;
        RECT 116.995 168.955 117.195 169.125 ;
        RECT 117.860 169.085 118.085 169.125 ;
        RECT 118.255 169.115 119.465 169.865 ;
        RECT 115.950 168.625 116.825 168.955 ;
        RECT 116.995 168.625 117.745 168.955 ;
        RECT 114.760 167.485 115.010 167.815 ;
        RECT 115.950 167.785 116.120 168.625 ;
        RECT 116.995 168.420 117.185 168.625 ;
        RECT 117.915 168.505 118.085 169.085 ;
        RECT 117.870 168.455 118.085 168.505 ;
        RECT 116.290 168.045 117.185 168.420 ;
        RECT 117.695 168.375 118.085 168.455 ;
        RECT 118.255 168.405 118.775 168.945 ;
        RECT 118.945 168.575 119.465 169.115 ;
        RECT 115.235 167.615 116.120 167.785 ;
        RECT 116.300 167.315 116.615 167.815 ;
        RECT 116.845 167.485 117.185 168.045 ;
        RECT 117.355 167.315 117.525 168.325 ;
        RECT 117.695 167.530 118.025 168.375 ;
        RECT 118.255 167.315 119.465 168.405 ;
        RECT 71.250 167.145 119.550 167.315 ;
        RECT 71.335 166.055 72.545 167.145 ;
        RECT 72.715 166.055 74.385 167.145 ;
        RECT 74.575 166.635 74.875 167.145 ;
        RECT 75.045 166.635 75.425 166.805 ;
        RECT 76.005 166.635 76.635 167.145 ;
        RECT 75.045 166.465 75.215 166.635 ;
        RECT 76.805 166.465 77.135 166.975 ;
        RECT 77.305 166.635 77.605 167.145 ;
        RECT 77.795 166.635 78.095 167.145 ;
        RECT 78.265 166.635 78.645 166.805 ;
        RECT 79.225 166.635 79.855 167.145 ;
        RECT 78.265 166.465 78.435 166.635 ;
        RECT 80.025 166.465 80.355 166.975 ;
        RECT 80.525 166.635 80.825 167.145 ;
        RECT 71.335 165.345 71.855 165.885 ;
        RECT 72.025 165.515 72.545 166.055 ;
        RECT 72.715 165.365 73.465 165.885 ;
        RECT 73.635 165.535 74.385 166.055 ;
        RECT 74.555 166.265 75.215 166.465 ;
        RECT 75.385 166.295 77.605 166.465 ;
        RECT 71.335 164.595 72.545 165.345 ;
        RECT 72.715 164.595 74.385 165.365 ;
        RECT 74.555 165.335 74.725 166.265 ;
        RECT 75.385 166.095 75.555 166.295 ;
        RECT 74.895 165.925 75.555 166.095 ;
        RECT 75.725 165.955 77.265 166.125 ;
        RECT 74.895 165.505 75.065 165.925 ;
        RECT 75.725 165.755 75.895 165.955 ;
        RECT 75.295 165.585 75.895 165.755 ;
        RECT 76.065 165.585 76.760 165.785 ;
        RECT 77.020 165.505 77.265 165.955 ;
        RECT 75.385 165.335 76.295 165.415 ;
        RECT 74.555 164.855 74.875 165.335 ;
        RECT 75.045 165.245 76.295 165.335 ;
        RECT 75.045 165.165 75.555 165.245 ;
        RECT 75.045 164.765 75.275 165.165 ;
        RECT 75.445 164.595 75.795 164.985 ;
        RECT 75.965 164.765 76.295 165.245 ;
        RECT 76.465 164.595 76.635 165.415 ;
        RECT 77.435 165.335 77.605 166.295 ;
        RECT 77.140 164.790 77.605 165.335 ;
        RECT 77.775 166.265 78.435 166.465 ;
        RECT 78.605 166.295 80.825 166.465 ;
        RECT 77.775 165.335 77.945 166.265 ;
        RECT 78.605 166.095 78.775 166.295 ;
        RECT 78.115 165.925 78.775 166.095 ;
        RECT 78.945 165.955 80.485 166.125 ;
        RECT 78.115 165.505 78.285 165.925 ;
        RECT 78.945 165.755 79.115 165.955 ;
        RECT 78.515 165.585 79.115 165.755 ;
        RECT 79.285 165.585 79.980 165.785 ;
        RECT 80.240 165.505 80.485 165.955 ;
        RECT 78.605 165.335 79.515 165.415 ;
        RECT 77.775 164.855 78.095 165.335 ;
        RECT 78.265 165.245 79.515 165.335 ;
        RECT 78.265 165.165 78.775 165.245 ;
        RECT 78.265 164.765 78.495 165.165 ;
        RECT 78.665 164.595 79.015 164.985 ;
        RECT 79.185 164.765 79.515 165.245 ;
        RECT 79.685 164.595 79.855 165.415 ;
        RECT 80.655 165.335 80.825 166.295 ;
        RECT 80.360 164.790 80.825 165.335 ;
        RECT 80.995 166.295 81.375 166.975 ;
        RECT 81.965 166.295 82.135 167.145 ;
        RECT 82.305 166.465 82.635 166.975 ;
        RECT 82.805 166.635 82.975 167.145 ;
        RECT 83.145 166.465 83.545 166.975 ;
        RECT 82.305 166.295 83.545 166.465 ;
        RECT 80.995 165.335 81.165 166.295 ;
        RECT 81.335 165.955 82.640 166.125 ;
        RECT 83.725 166.045 84.045 166.975 ;
        RECT 81.335 165.505 81.580 165.955 ;
        RECT 81.750 165.585 82.300 165.785 ;
        RECT 82.470 165.755 82.640 165.955 ;
        RECT 83.415 165.875 84.045 166.045 ;
        RECT 84.215 165.980 84.505 167.145 ;
        RECT 84.675 166.055 85.885 167.145 ;
        RECT 86.170 166.515 86.455 166.975 ;
        RECT 86.625 166.685 86.895 167.145 ;
        RECT 86.170 166.295 87.125 166.515 ;
        RECT 82.470 165.585 82.845 165.755 ;
        RECT 83.015 165.335 83.245 165.835 ;
        RECT 80.995 165.165 83.245 165.335 ;
        RECT 81.045 164.595 81.375 164.985 ;
        RECT 81.545 164.845 81.715 165.165 ;
        RECT 83.415 164.995 83.585 165.875 ;
        RECT 81.885 164.595 82.215 164.985 ;
        RECT 82.630 164.825 83.585 164.995 ;
        RECT 83.755 164.595 84.045 165.430 ;
        RECT 84.675 165.345 85.195 165.885 ;
        RECT 85.365 165.515 85.885 166.055 ;
        RECT 86.055 165.565 86.745 166.125 ;
        RECT 86.915 165.395 87.125 166.295 ;
        RECT 84.215 164.595 84.505 165.320 ;
        RECT 84.675 164.595 85.885 165.345 ;
        RECT 86.170 165.225 87.125 165.395 ;
        RECT 87.295 166.125 87.695 166.975 ;
        RECT 87.885 166.515 88.165 166.975 ;
        RECT 88.685 166.685 89.010 167.145 ;
        RECT 87.885 166.295 89.010 166.515 ;
        RECT 87.295 165.565 88.390 166.125 ;
        RECT 88.560 165.835 89.010 166.295 ;
        RECT 89.180 166.005 89.565 166.975 ;
        RECT 89.735 166.055 91.405 167.145 ;
        RECT 86.170 164.765 86.455 165.225 ;
        RECT 86.625 164.595 86.895 165.055 ;
        RECT 87.295 164.765 87.695 165.565 ;
        RECT 88.560 165.505 89.115 165.835 ;
        RECT 88.560 165.395 89.010 165.505 ;
        RECT 87.885 165.225 89.010 165.395 ;
        RECT 89.285 165.335 89.565 166.005 ;
        RECT 87.885 164.765 88.165 165.225 ;
        RECT 88.685 164.595 89.010 165.055 ;
        RECT 89.180 164.765 89.565 165.335 ;
        RECT 89.735 165.365 90.485 165.885 ;
        RECT 90.655 165.535 91.405 166.055 ;
        RECT 92.035 166.070 92.305 166.975 ;
        RECT 92.475 166.385 92.805 167.145 ;
        RECT 92.985 166.215 93.165 166.975 ;
        RECT 93.420 166.475 93.675 166.975 ;
        RECT 93.845 166.645 94.175 167.145 ;
        RECT 93.420 166.305 94.170 166.475 ;
        RECT 89.735 164.595 91.405 165.365 ;
        RECT 92.035 165.270 92.215 166.070 ;
        RECT 92.490 166.045 93.165 166.215 ;
        RECT 92.490 165.900 92.660 166.045 ;
        RECT 92.385 165.570 92.660 165.900 ;
        RECT 92.490 165.315 92.660 165.570 ;
        RECT 92.885 165.495 93.225 165.865 ;
        RECT 93.420 165.485 93.770 166.135 ;
        RECT 93.940 165.315 94.170 166.305 ;
        RECT 92.035 164.765 92.295 165.270 ;
        RECT 92.490 165.145 93.155 165.315 ;
        RECT 92.475 164.595 92.805 164.975 ;
        RECT 92.985 164.765 93.155 165.145 ;
        RECT 93.420 165.145 94.170 165.315 ;
        RECT 93.420 164.855 93.675 165.145 ;
        RECT 93.845 164.595 94.175 164.975 ;
        RECT 94.345 164.855 94.515 166.975 ;
        RECT 94.685 166.175 95.010 166.960 ;
        RECT 95.180 166.685 95.430 167.145 ;
        RECT 95.600 166.645 95.850 166.975 ;
        RECT 96.065 166.645 96.745 166.975 ;
        RECT 95.600 166.515 95.770 166.645 ;
        RECT 95.375 166.345 95.770 166.515 ;
        RECT 94.745 165.125 95.205 166.175 ;
        RECT 95.375 164.985 95.545 166.345 ;
        RECT 95.940 166.085 96.405 166.475 ;
        RECT 95.715 165.275 96.065 165.895 ;
        RECT 96.235 165.495 96.405 166.085 ;
        RECT 96.575 165.865 96.745 166.645 ;
        RECT 96.915 166.545 97.085 166.885 ;
        RECT 97.320 166.715 97.650 167.145 ;
        RECT 97.820 166.545 97.990 166.885 ;
        RECT 98.285 166.685 98.655 167.145 ;
        RECT 96.915 166.375 97.990 166.545 ;
        RECT 98.825 166.515 98.995 166.975 ;
        RECT 99.230 166.635 100.100 166.975 ;
        RECT 100.270 166.685 100.520 167.145 ;
        RECT 98.435 166.345 98.995 166.515 ;
        RECT 98.435 166.205 98.605 166.345 ;
        RECT 97.105 166.035 98.605 166.205 ;
        RECT 99.300 166.175 99.760 166.465 ;
        RECT 96.575 165.695 98.265 165.865 ;
        RECT 96.235 165.275 96.590 165.495 ;
        RECT 96.760 164.985 96.930 165.695 ;
        RECT 97.135 165.275 97.925 165.525 ;
        RECT 98.095 165.515 98.265 165.695 ;
        RECT 98.435 165.345 98.605 166.035 ;
        RECT 94.875 164.595 95.205 164.955 ;
        RECT 95.375 164.815 95.870 164.985 ;
        RECT 96.075 164.815 96.930 164.985 ;
        RECT 97.805 164.595 98.135 165.055 ;
        RECT 98.345 164.955 98.605 165.345 ;
        RECT 98.795 166.165 99.760 166.175 ;
        RECT 99.930 166.255 100.100 166.635 ;
        RECT 100.690 166.595 100.860 166.885 ;
        RECT 101.040 166.765 101.370 167.145 ;
        RECT 100.690 166.425 101.490 166.595 ;
        RECT 98.795 166.005 99.470 166.165 ;
        RECT 99.930 166.085 101.150 166.255 ;
        RECT 98.795 165.215 99.005 166.005 ;
        RECT 99.930 165.995 100.100 166.085 ;
        RECT 99.175 165.215 99.525 165.835 ;
        RECT 99.695 165.825 100.100 165.995 ;
        RECT 99.695 165.045 99.865 165.825 ;
        RECT 100.035 165.375 100.255 165.655 ;
        RECT 100.435 165.545 100.975 165.915 ;
        RECT 101.320 165.835 101.490 166.425 ;
        RECT 101.710 166.005 102.015 167.145 ;
        RECT 102.185 165.955 102.440 166.835 ;
        RECT 102.615 166.055 106.125 167.145 ;
        RECT 101.320 165.805 102.060 165.835 ;
        RECT 100.035 165.205 100.565 165.375 ;
        RECT 98.345 164.785 98.695 164.955 ;
        RECT 98.915 164.765 99.865 165.045 ;
        RECT 100.035 164.595 100.225 165.035 ;
        RECT 100.395 164.975 100.565 165.205 ;
        RECT 100.735 165.145 100.975 165.545 ;
        RECT 101.145 165.505 102.060 165.805 ;
        RECT 101.145 165.330 101.470 165.505 ;
        RECT 101.145 164.975 101.465 165.330 ;
        RECT 102.230 165.305 102.440 165.955 ;
        RECT 100.395 164.805 101.465 164.975 ;
        RECT 101.710 164.595 102.015 165.055 ;
        RECT 102.185 164.775 102.440 165.305 ;
        RECT 102.615 165.365 104.265 165.885 ;
        RECT 104.435 165.535 106.125 166.055 ;
        RECT 106.755 166.005 107.025 166.975 ;
        RECT 107.235 166.345 107.515 167.145 ;
        RECT 107.695 166.595 108.890 166.925 ;
        RECT 108.020 166.175 108.440 166.425 ;
        RECT 107.195 166.005 108.440 166.175 ;
        RECT 102.615 164.595 106.125 165.365 ;
        RECT 106.755 165.270 106.925 166.005 ;
        RECT 107.195 165.835 107.365 166.005 ;
        RECT 108.665 165.835 108.835 166.395 ;
        RECT 109.085 166.005 109.340 167.145 ;
        RECT 109.975 165.980 110.265 167.145 ;
        RECT 110.435 166.055 111.645 167.145 ;
        RECT 107.135 165.505 107.365 165.835 ;
        RECT 108.095 165.505 108.835 165.835 ;
        RECT 109.005 165.585 109.340 165.835 ;
        RECT 107.195 165.335 107.365 165.505 ;
        RECT 108.585 165.415 108.835 165.505 ;
        RECT 106.755 164.925 107.025 165.270 ;
        RECT 107.195 165.165 107.935 165.335 ;
        RECT 108.585 165.245 109.320 165.415 ;
        RECT 110.435 165.345 110.955 165.885 ;
        RECT 111.125 165.515 111.645 166.055 ;
        RECT 111.815 166.005 112.200 166.975 ;
        RECT 112.370 166.685 112.695 167.145 ;
        RECT 113.215 166.515 113.495 166.975 ;
        RECT 112.370 166.295 113.495 166.515 ;
        RECT 107.215 164.595 107.595 164.995 ;
        RECT 107.765 164.815 107.935 165.165 ;
        RECT 108.105 164.595 108.840 165.075 ;
        RECT 109.010 164.775 109.320 165.245 ;
        RECT 109.975 164.595 110.265 165.320 ;
        RECT 110.435 164.595 111.645 165.345 ;
        RECT 111.815 165.335 112.095 166.005 ;
        RECT 112.370 165.835 112.820 166.295 ;
        RECT 113.685 166.125 114.085 166.975 ;
        RECT 114.485 166.685 114.755 167.145 ;
        RECT 114.925 166.515 115.210 166.975 ;
        RECT 112.265 165.505 112.820 165.835 ;
        RECT 112.990 165.565 114.085 166.125 ;
        RECT 112.370 165.395 112.820 165.505 ;
        RECT 111.815 164.765 112.200 165.335 ;
        RECT 112.370 165.225 113.495 165.395 ;
        RECT 112.370 164.595 112.695 165.055 ;
        RECT 113.215 164.765 113.495 165.225 ;
        RECT 113.685 164.765 114.085 165.565 ;
        RECT 114.255 166.295 115.210 166.515 ;
        RECT 114.255 165.395 114.465 166.295 ;
        RECT 114.635 165.565 115.325 166.125 ;
        RECT 115.495 166.005 115.755 167.145 ;
        RECT 115.925 165.995 116.255 166.975 ;
        RECT 116.425 166.005 116.705 167.145 ;
        RECT 116.875 166.055 118.085 167.145 ;
        RECT 115.515 165.585 115.850 165.835 ;
        RECT 116.020 165.395 116.190 165.995 ;
        RECT 116.360 165.565 116.695 165.835 ;
        RECT 114.255 165.225 115.210 165.395 ;
        RECT 114.485 164.595 114.755 165.055 ;
        RECT 114.925 164.765 115.210 165.225 ;
        RECT 115.495 164.765 116.190 165.395 ;
        RECT 116.395 164.595 116.705 165.395 ;
        RECT 116.875 165.345 117.395 165.885 ;
        RECT 117.565 165.515 118.085 166.055 ;
        RECT 118.255 166.055 119.465 167.145 ;
        RECT 118.255 165.515 118.775 166.055 ;
        RECT 118.945 165.345 119.465 165.885 ;
        RECT 116.875 164.595 118.085 165.345 ;
        RECT 118.255 164.595 119.465 165.345 ;
        RECT 71.250 164.425 119.550 164.595 ;
        RECT 71.335 163.675 72.545 164.425 ;
        RECT 71.335 163.135 71.855 163.675 ;
        RECT 72.715 163.655 75.305 164.425 ;
        RECT 75.480 163.875 75.735 164.165 ;
        RECT 75.905 164.045 76.235 164.425 ;
        RECT 75.480 163.705 76.230 163.875 ;
        RECT 72.025 162.965 72.545 163.505 ;
        RECT 72.715 163.135 73.925 163.655 ;
        RECT 74.095 162.965 75.305 163.485 ;
        RECT 71.335 161.875 72.545 162.965 ;
        RECT 72.715 161.875 75.305 162.965 ;
        RECT 75.480 162.885 75.830 163.535 ;
        RECT 76.000 162.715 76.230 163.705 ;
        RECT 75.480 162.545 76.230 162.715 ;
        RECT 75.480 162.045 75.735 162.545 ;
        RECT 75.905 161.875 76.235 162.375 ;
        RECT 76.405 162.045 76.575 164.165 ;
        RECT 76.935 164.065 77.265 164.425 ;
        RECT 77.435 164.035 77.930 164.205 ;
        RECT 78.135 164.035 78.990 164.205 ;
        RECT 76.805 162.845 77.265 163.895 ;
        RECT 76.745 162.060 77.070 162.845 ;
        RECT 77.435 162.675 77.605 164.035 ;
        RECT 77.775 163.125 78.125 163.745 ;
        RECT 78.295 163.525 78.650 163.745 ;
        RECT 78.295 162.935 78.465 163.525 ;
        RECT 78.820 163.325 78.990 164.035 ;
        RECT 79.865 163.965 80.195 164.425 ;
        RECT 80.405 164.065 80.755 164.235 ;
        RECT 79.195 163.495 79.985 163.745 ;
        RECT 80.405 163.675 80.665 164.065 ;
        RECT 80.975 163.975 81.925 164.255 ;
        RECT 82.095 163.985 82.285 164.425 ;
        RECT 82.455 164.045 83.525 164.215 ;
        RECT 80.155 163.325 80.325 163.505 ;
        RECT 77.435 162.505 77.830 162.675 ;
        RECT 78.000 162.545 78.465 162.935 ;
        RECT 78.635 163.155 80.325 163.325 ;
        RECT 77.660 162.375 77.830 162.505 ;
        RECT 78.635 162.375 78.805 163.155 ;
        RECT 80.495 162.985 80.665 163.675 ;
        RECT 79.165 162.815 80.665 162.985 ;
        RECT 80.855 163.015 81.065 163.805 ;
        RECT 81.235 163.185 81.585 163.805 ;
        RECT 81.755 163.195 81.925 163.975 ;
        RECT 82.455 163.815 82.625 164.045 ;
        RECT 82.095 163.645 82.625 163.815 ;
        RECT 82.095 163.365 82.315 163.645 ;
        RECT 82.795 163.475 83.035 163.875 ;
        RECT 81.755 163.025 82.160 163.195 ;
        RECT 82.495 163.105 83.035 163.475 ;
        RECT 83.205 163.690 83.525 164.045 ;
        RECT 83.770 163.965 84.075 164.425 ;
        RECT 84.245 163.715 84.500 164.245 ;
        RECT 83.205 163.515 83.530 163.690 ;
        RECT 83.205 163.215 84.120 163.515 ;
        RECT 83.380 163.185 84.120 163.215 ;
        RECT 80.855 162.855 81.530 163.015 ;
        RECT 81.990 162.935 82.160 163.025 ;
        RECT 80.855 162.845 81.820 162.855 ;
        RECT 80.495 162.675 80.665 162.815 ;
        RECT 77.240 161.875 77.490 162.335 ;
        RECT 77.660 162.045 77.910 162.375 ;
        RECT 78.125 162.045 78.805 162.375 ;
        RECT 78.975 162.475 80.050 162.645 ;
        RECT 80.495 162.505 81.055 162.675 ;
        RECT 81.360 162.555 81.820 162.845 ;
        RECT 81.990 162.765 83.210 162.935 ;
        RECT 78.975 162.135 79.145 162.475 ;
        RECT 79.380 161.875 79.710 162.305 ;
        RECT 79.880 162.135 80.050 162.475 ;
        RECT 80.345 161.875 80.715 162.335 ;
        RECT 80.885 162.045 81.055 162.505 ;
        RECT 81.990 162.385 82.160 162.765 ;
        RECT 83.380 162.595 83.550 163.185 ;
        RECT 84.290 163.065 84.500 163.715 ;
        RECT 81.290 162.045 82.160 162.385 ;
        RECT 82.750 162.425 83.550 162.595 ;
        RECT 82.330 161.875 82.580 162.335 ;
        RECT 82.750 162.135 82.920 162.425 ;
        RECT 83.100 161.875 83.430 162.255 ;
        RECT 83.770 161.875 84.075 163.015 ;
        RECT 84.245 162.185 84.500 163.065 ;
        RECT 85.600 163.715 85.855 164.245 ;
        RECT 86.025 163.965 86.330 164.425 ;
        RECT 86.575 164.045 87.645 164.215 ;
        RECT 85.600 163.065 85.810 163.715 ;
        RECT 86.575 163.690 86.895 164.045 ;
        RECT 86.570 163.515 86.895 163.690 ;
        RECT 85.980 163.215 86.895 163.515 ;
        RECT 87.065 163.475 87.305 163.875 ;
        RECT 87.475 163.815 87.645 164.045 ;
        RECT 87.815 163.985 88.005 164.425 ;
        RECT 88.175 163.975 89.125 164.255 ;
        RECT 89.345 164.065 89.695 164.235 ;
        RECT 87.475 163.645 88.005 163.815 ;
        RECT 85.980 163.185 86.720 163.215 ;
        RECT 85.600 162.185 85.855 163.065 ;
        RECT 86.025 161.875 86.330 163.015 ;
        RECT 86.550 162.595 86.720 163.185 ;
        RECT 87.065 163.105 87.605 163.475 ;
        RECT 87.785 163.365 88.005 163.645 ;
        RECT 88.175 163.195 88.345 163.975 ;
        RECT 87.940 163.025 88.345 163.195 ;
        RECT 88.515 163.185 88.865 163.805 ;
        RECT 87.940 162.935 88.110 163.025 ;
        RECT 89.035 163.015 89.245 163.805 ;
        RECT 86.890 162.765 88.110 162.935 ;
        RECT 88.570 162.855 89.245 163.015 ;
        RECT 86.550 162.425 87.350 162.595 ;
        RECT 86.670 161.875 87.000 162.255 ;
        RECT 87.180 162.135 87.350 162.425 ;
        RECT 87.940 162.385 88.110 162.765 ;
        RECT 88.280 162.845 89.245 162.855 ;
        RECT 89.435 163.675 89.695 164.065 ;
        RECT 89.905 163.965 90.235 164.425 ;
        RECT 91.110 164.035 91.965 164.205 ;
        RECT 92.170 164.035 92.665 164.205 ;
        RECT 92.835 164.065 93.165 164.425 ;
        RECT 89.435 162.985 89.605 163.675 ;
        RECT 89.775 163.325 89.945 163.505 ;
        RECT 90.115 163.495 90.905 163.745 ;
        RECT 91.110 163.325 91.280 164.035 ;
        RECT 91.450 163.525 91.805 163.745 ;
        RECT 89.775 163.155 91.465 163.325 ;
        RECT 88.280 162.555 88.740 162.845 ;
        RECT 89.435 162.815 90.935 162.985 ;
        RECT 89.435 162.675 89.605 162.815 ;
        RECT 89.045 162.505 89.605 162.675 ;
        RECT 87.520 161.875 87.770 162.335 ;
        RECT 87.940 162.045 88.810 162.385 ;
        RECT 89.045 162.045 89.215 162.505 ;
        RECT 90.050 162.475 91.125 162.645 ;
        RECT 89.385 161.875 89.755 162.335 ;
        RECT 90.050 162.135 90.220 162.475 ;
        RECT 90.390 161.875 90.720 162.305 ;
        RECT 90.955 162.135 91.125 162.475 ;
        RECT 91.295 162.375 91.465 163.155 ;
        RECT 91.635 162.935 91.805 163.525 ;
        RECT 91.975 163.125 92.325 163.745 ;
        RECT 91.635 162.545 92.100 162.935 ;
        RECT 92.495 162.675 92.665 164.035 ;
        RECT 92.835 162.845 93.295 163.895 ;
        RECT 92.270 162.505 92.665 162.675 ;
        RECT 92.270 162.375 92.440 162.505 ;
        RECT 91.295 162.045 91.975 162.375 ;
        RECT 92.190 162.045 92.440 162.375 ;
        RECT 92.610 161.875 92.860 162.335 ;
        RECT 93.030 162.060 93.355 162.845 ;
        RECT 93.525 162.045 93.695 164.165 ;
        RECT 93.865 164.045 94.195 164.425 ;
        RECT 94.365 163.875 94.620 164.165 ;
        RECT 93.870 163.705 94.620 163.875 ;
        RECT 93.870 162.715 94.100 163.705 ;
        RECT 94.795 163.655 96.465 164.425 ;
        RECT 97.095 163.700 97.385 164.425 ;
        RECT 97.560 163.875 97.815 164.165 ;
        RECT 97.985 164.045 98.315 164.425 ;
        RECT 97.560 163.705 98.310 163.875 ;
        RECT 94.270 162.885 94.620 163.535 ;
        RECT 94.795 163.135 95.545 163.655 ;
        RECT 95.715 162.965 96.465 163.485 ;
        RECT 93.870 162.545 94.620 162.715 ;
        RECT 93.865 161.875 94.195 162.375 ;
        RECT 94.365 162.045 94.620 162.545 ;
        RECT 94.795 161.875 96.465 162.965 ;
        RECT 97.095 161.875 97.385 163.040 ;
        RECT 97.560 162.885 97.910 163.535 ;
        RECT 98.080 162.715 98.310 163.705 ;
        RECT 97.560 162.545 98.310 162.715 ;
        RECT 97.560 162.045 97.815 162.545 ;
        RECT 97.985 161.875 98.315 162.375 ;
        RECT 98.485 162.045 98.655 164.165 ;
        RECT 99.015 164.065 99.345 164.425 ;
        RECT 99.515 164.035 100.010 164.205 ;
        RECT 100.215 164.035 101.070 164.205 ;
        RECT 98.885 162.845 99.345 163.895 ;
        RECT 98.825 162.060 99.150 162.845 ;
        RECT 99.515 162.675 99.685 164.035 ;
        RECT 99.855 163.125 100.205 163.745 ;
        RECT 100.375 163.525 100.730 163.745 ;
        RECT 100.375 162.935 100.545 163.525 ;
        RECT 100.900 163.325 101.070 164.035 ;
        RECT 101.945 163.965 102.275 164.425 ;
        RECT 102.485 164.065 102.835 164.235 ;
        RECT 101.275 163.495 102.065 163.745 ;
        RECT 102.485 163.675 102.745 164.065 ;
        RECT 103.055 163.975 104.005 164.255 ;
        RECT 104.175 163.985 104.365 164.425 ;
        RECT 104.535 164.045 105.605 164.215 ;
        RECT 102.235 163.325 102.405 163.505 ;
        RECT 99.515 162.505 99.910 162.675 ;
        RECT 100.080 162.545 100.545 162.935 ;
        RECT 100.715 163.155 102.405 163.325 ;
        RECT 99.740 162.375 99.910 162.505 ;
        RECT 100.715 162.375 100.885 163.155 ;
        RECT 102.575 162.985 102.745 163.675 ;
        RECT 101.245 162.815 102.745 162.985 ;
        RECT 102.935 163.015 103.145 163.805 ;
        RECT 103.315 163.185 103.665 163.805 ;
        RECT 103.835 163.195 104.005 163.975 ;
        RECT 104.535 163.815 104.705 164.045 ;
        RECT 104.175 163.645 104.705 163.815 ;
        RECT 104.175 163.365 104.395 163.645 ;
        RECT 104.875 163.475 105.115 163.875 ;
        RECT 103.835 163.025 104.240 163.195 ;
        RECT 104.575 163.105 105.115 163.475 ;
        RECT 105.285 163.690 105.605 164.045 ;
        RECT 105.850 163.965 106.155 164.425 ;
        RECT 106.325 163.715 106.580 164.245 ;
        RECT 105.285 163.515 105.610 163.690 ;
        RECT 105.285 163.215 106.200 163.515 ;
        RECT 105.460 163.185 106.200 163.215 ;
        RECT 102.935 162.855 103.610 163.015 ;
        RECT 104.070 162.935 104.240 163.025 ;
        RECT 102.935 162.845 103.900 162.855 ;
        RECT 102.575 162.675 102.745 162.815 ;
        RECT 99.320 161.875 99.570 162.335 ;
        RECT 99.740 162.045 99.990 162.375 ;
        RECT 100.205 162.045 100.885 162.375 ;
        RECT 101.055 162.475 102.130 162.645 ;
        RECT 102.575 162.505 103.135 162.675 ;
        RECT 103.440 162.555 103.900 162.845 ;
        RECT 104.070 162.765 105.290 162.935 ;
        RECT 101.055 162.135 101.225 162.475 ;
        RECT 101.460 161.875 101.790 162.305 ;
        RECT 101.960 162.135 102.130 162.475 ;
        RECT 102.425 161.875 102.795 162.335 ;
        RECT 102.965 162.045 103.135 162.505 ;
        RECT 104.070 162.385 104.240 162.765 ;
        RECT 105.460 162.595 105.630 163.185 ;
        RECT 106.370 163.065 106.580 163.715 ;
        RECT 106.755 163.675 107.965 164.425 ;
        RECT 108.225 163.875 108.395 164.165 ;
        RECT 108.565 164.045 108.895 164.425 ;
        RECT 108.225 163.705 108.890 163.875 ;
        RECT 106.755 163.135 107.275 163.675 ;
        RECT 103.370 162.045 104.240 162.385 ;
        RECT 104.830 162.425 105.630 162.595 ;
        RECT 104.410 161.875 104.660 162.335 ;
        RECT 104.830 162.135 105.000 162.425 ;
        RECT 105.180 161.875 105.510 162.255 ;
        RECT 105.850 161.875 106.155 163.015 ;
        RECT 106.325 162.185 106.580 163.065 ;
        RECT 107.445 162.965 107.965 163.505 ;
        RECT 106.755 161.875 107.965 162.965 ;
        RECT 108.140 162.885 108.490 163.535 ;
        RECT 108.660 162.715 108.890 163.705 ;
        RECT 108.225 162.545 108.890 162.715 ;
        RECT 108.225 162.045 108.395 162.545 ;
        RECT 108.565 161.875 108.895 162.375 ;
        RECT 109.065 162.045 109.250 164.165 ;
        RECT 109.505 163.965 109.755 164.425 ;
        RECT 109.925 163.975 110.260 164.145 ;
        RECT 110.455 163.975 111.130 164.145 ;
        RECT 109.925 163.835 110.095 163.975 ;
        RECT 109.420 162.845 109.700 163.795 ;
        RECT 109.870 163.705 110.095 163.835 ;
        RECT 109.870 162.600 110.040 163.705 ;
        RECT 110.265 163.555 110.790 163.775 ;
        RECT 110.210 162.790 110.450 163.385 ;
        RECT 110.620 162.855 110.790 163.555 ;
        RECT 110.960 163.195 111.130 163.975 ;
        RECT 111.450 163.925 111.820 164.425 ;
        RECT 112.000 163.975 112.405 164.145 ;
        RECT 112.575 163.975 113.360 164.145 ;
        RECT 112.000 163.745 112.170 163.975 ;
        RECT 111.340 163.445 112.170 163.745 ;
        RECT 112.555 163.475 113.020 163.805 ;
        RECT 111.340 163.415 111.540 163.445 ;
        RECT 111.660 163.195 111.830 163.265 ;
        RECT 110.960 163.025 111.830 163.195 ;
        RECT 111.320 162.935 111.830 163.025 ;
        RECT 109.870 162.470 110.175 162.600 ;
        RECT 110.620 162.490 111.150 162.855 ;
        RECT 109.490 161.875 109.755 162.335 ;
        RECT 109.925 162.045 110.175 162.470 ;
        RECT 111.320 162.320 111.490 162.935 ;
        RECT 110.385 162.150 111.490 162.320 ;
        RECT 111.660 161.875 111.830 162.675 ;
        RECT 112.000 162.375 112.170 163.445 ;
        RECT 112.340 162.545 112.530 163.265 ;
        RECT 112.700 162.515 113.020 163.475 ;
        RECT 113.190 163.515 113.360 163.975 ;
        RECT 113.635 163.895 113.845 164.425 ;
        RECT 114.105 163.685 114.435 164.210 ;
        RECT 114.605 163.815 114.775 164.425 ;
        RECT 114.945 163.770 115.275 164.205 ;
        RECT 114.945 163.685 115.325 163.770 ;
        RECT 114.235 163.515 114.435 163.685 ;
        RECT 115.100 163.645 115.325 163.685 ;
        RECT 113.190 163.185 114.065 163.515 ;
        RECT 114.235 163.185 114.985 163.515 ;
        RECT 112.000 162.045 112.250 162.375 ;
        RECT 113.190 162.345 113.360 163.185 ;
        RECT 114.235 162.980 114.425 163.185 ;
        RECT 115.155 163.065 115.325 163.645 ;
        RECT 115.495 163.655 118.085 164.425 ;
        RECT 118.255 163.675 119.465 164.425 ;
        RECT 115.495 163.135 116.705 163.655 ;
        RECT 115.110 163.015 115.325 163.065 ;
        RECT 113.530 162.605 114.425 162.980 ;
        RECT 114.935 162.935 115.325 163.015 ;
        RECT 116.875 162.965 118.085 163.485 ;
        RECT 112.475 162.175 113.360 162.345 ;
        RECT 113.540 161.875 113.855 162.375 ;
        RECT 114.085 162.045 114.425 162.605 ;
        RECT 114.595 161.875 114.765 162.885 ;
        RECT 114.935 162.090 115.265 162.935 ;
        RECT 115.495 161.875 118.085 162.965 ;
        RECT 118.255 162.965 118.775 163.505 ;
        RECT 118.945 163.135 119.465 163.675 ;
        RECT 118.255 161.875 119.465 162.965 ;
        RECT 71.250 161.705 119.550 161.875 ;
        RECT 71.335 160.615 72.545 161.705 ;
        RECT 72.715 161.270 78.060 161.705 ;
        RECT 78.235 161.270 83.580 161.705 ;
        RECT 71.335 159.905 71.855 160.445 ;
        RECT 72.025 160.075 72.545 160.615 ;
        RECT 71.335 159.155 72.545 159.905 ;
        RECT 74.300 159.700 74.640 160.530 ;
        RECT 76.120 160.020 76.470 161.270 ;
        RECT 79.820 159.700 80.160 160.530 ;
        RECT 81.640 160.020 81.990 161.270 ;
        RECT 84.215 160.540 84.505 161.705 ;
        RECT 84.675 160.615 86.345 161.705 ;
        RECT 86.515 161.110 86.950 161.535 ;
        RECT 87.120 161.280 87.505 161.705 ;
        RECT 86.515 160.940 87.505 161.110 ;
        RECT 84.675 159.925 85.425 160.445 ;
        RECT 85.595 160.095 86.345 160.615 ;
        RECT 86.515 160.065 87.000 160.770 ;
        RECT 87.170 160.395 87.505 160.940 ;
        RECT 87.675 160.745 88.100 161.535 ;
        RECT 88.270 161.110 88.545 161.535 ;
        RECT 88.715 161.280 89.100 161.705 ;
        RECT 88.270 160.915 89.100 161.110 ;
        RECT 87.675 160.565 88.580 160.745 ;
        RECT 87.170 160.065 87.580 160.395 ;
        RECT 87.750 160.065 88.580 160.565 ;
        RECT 88.750 160.395 89.100 160.915 ;
        RECT 89.270 160.745 89.515 161.535 ;
        RECT 89.705 161.110 89.960 161.535 ;
        RECT 90.130 161.280 90.515 161.705 ;
        RECT 89.705 160.915 90.515 161.110 ;
        RECT 89.270 160.565 89.995 160.745 ;
        RECT 88.750 160.065 89.175 160.395 ;
        RECT 89.345 160.065 89.995 160.565 ;
        RECT 90.165 160.395 90.515 160.915 ;
        RECT 90.685 160.565 90.945 161.535 ;
        RECT 91.115 161.270 96.460 161.705 ;
        RECT 96.635 161.270 101.980 161.705 ;
        RECT 90.165 160.065 90.590 160.395 ;
        RECT 72.715 159.155 78.060 159.700 ;
        RECT 78.235 159.155 83.580 159.700 ;
        RECT 84.215 159.155 84.505 159.880 ;
        RECT 84.675 159.155 86.345 159.925 ;
        RECT 87.170 159.895 87.505 160.065 ;
        RECT 87.750 159.895 88.100 160.065 ;
        RECT 88.750 159.895 89.100 160.065 ;
        RECT 89.345 159.895 89.515 160.065 ;
        RECT 90.165 159.895 90.515 160.065 ;
        RECT 90.760 159.895 90.945 160.565 ;
        RECT 86.515 159.725 87.505 159.895 ;
        RECT 86.515 159.325 86.950 159.725 ;
        RECT 87.120 159.155 87.505 159.555 ;
        RECT 87.675 159.325 88.100 159.895 ;
        RECT 88.290 159.725 89.100 159.895 ;
        RECT 88.290 159.325 88.545 159.725 ;
        RECT 88.715 159.155 89.100 159.555 ;
        RECT 89.270 159.325 89.515 159.895 ;
        RECT 89.705 159.725 90.515 159.895 ;
        RECT 89.705 159.325 89.960 159.725 ;
        RECT 90.130 159.155 90.515 159.555 ;
        RECT 90.685 159.325 90.945 159.895 ;
        RECT 92.700 159.700 93.040 160.530 ;
        RECT 94.520 160.020 94.870 161.270 ;
        RECT 98.220 159.700 98.560 160.530 ;
        RECT 100.040 160.020 100.390 161.270 ;
        RECT 102.270 161.075 102.555 161.535 ;
        RECT 102.725 161.245 102.995 161.705 ;
        RECT 102.270 160.855 103.225 161.075 ;
        RECT 102.155 160.125 102.845 160.685 ;
        RECT 103.015 159.955 103.225 160.855 ;
        RECT 102.270 159.785 103.225 159.955 ;
        RECT 103.395 160.685 103.795 161.535 ;
        RECT 103.985 161.075 104.265 161.535 ;
        RECT 104.785 161.245 105.110 161.705 ;
        RECT 103.985 160.855 105.110 161.075 ;
        RECT 103.395 160.125 104.490 160.685 ;
        RECT 104.660 160.395 105.110 160.855 ;
        RECT 105.280 160.565 105.665 161.535 ;
        RECT 91.115 159.155 96.460 159.700 ;
        RECT 96.635 159.155 101.980 159.700 ;
        RECT 102.270 159.325 102.555 159.785 ;
        RECT 102.725 159.155 102.995 159.615 ;
        RECT 103.395 159.325 103.795 160.125 ;
        RECT 104.660 160.065 105.215 160.395 ;
        RECT 104.660 159.955 105.110 160.065 ;
        RECT 103.985 159.785 105.110 159.955 ;
        RECT 105.385 159.895 105.665 160.565 ;
        RECT 103.985 159.325 104.265 159.785 ;
        RECT 104.785 159.155 105.110 159.615 ;
        RECT 105.280 159.325 105.665 159.895 ;
        RECT 105.835 160.565 106.220 161.535 ;
        RECT 106.390 161.245 106.715 161.705 ;
        RECT 107.235 161.075 107.515 161.535 ;
        RECT 106.390 160.855 107.515 161.075 ;
        RECT 105.835 159.895 106.115 160.565 ;
        RECT 106.390 160.395 106.840 160.855 ;
        RECT 107.705 160.685 108.105 161.535 ;
        RECT 108.505 161.245 108.775 161.705 ;
        RECT 108.945 161.075 109.230 161.535 ;
        RECT 106.285 160.065 106.840 160.395 ;
        RECT 107.010 160.125 108.105 160.685 ;
        RECT 106.390 159.955 106.840 160.065 ;
        RECT 105.835 159.325 106.220 159.895 ;
        RECT 106.390 159.785 107.515 159.955 ;
        RECT 106.390 159.155 106.715 159.615 ;
        RECT 107.235 159.325 107.515 159.785 ;
        RECT 107.705 159.325 108.105 160.125 ;
        RECT 108.275 160.855 109.230 161.075 ;
        RECT 108.275 159.955 108.485 160.855 ;
        RECT 108.655 160.125 109.345 160.685 ;
        RECT 109.975 160.540 110.265 161.705 ;
        RECT 110.555 160.585 110.885 161.705 ;
        RECT 110.495 160.145 111.005 160.395 ;
        RECT 111.215 160.145 111.585 161.460 ;
        RECT 111.755 160.145 112.085 161.460 ;
        RECT 112.295 160.145 112.625 161.460 ;
        RECT 112.895 160.815 113.145 161.535 ;
        RECT 113.315 160.985 113.645 161.705 ;
        RECT 112.895 160.525 113.645 160.815 ;
        RECT 113.880 160.525 114.405 161.535 ;
        RECT 113.385 160.355 113.645 160.525 ;
        RECT 112.795 160.145 113.215 160.355 ;
        RECT 113.385 160.145 113.965 160.355 ;
        RECT 113.385 159.975 113.755 160.145 ;
        RECT 108.275 159.785 109.230 159.955 ;
        RECT 108.505 159.155 108.775 159.615 ;
        RECT 108.945 159.325 109.230 159.785 ;
        RECT 109.975 159.155 110.265 159.880 ;
        RECT 110.535 159.805 112.835 159.975 ;
        RECT 110.535 159.325 110.865 159.805 ;
        RECT 111.035 159.155 111.365 159.615 ;
        RECT 111.580 159.325 111.910 159.805 ;
        RECT 112.110 159.155 112.440 159.615 ;
        RECT 112.665 159.485 112.835 159.805 ;
        RECT 113.005 159.785 113.755 159.975 ;
        RECT 114.135 159.955 114.405 160.525 ;
        RECT 113.005 159.340 113.335 159.785 ;
        RECT 113.605 159.155 113.775 159.615 ;
        RECT 114.065 159.325 114.405 159.955 ;
        RECT 114.575 160.565 114.960 161.535 ;
        RECT 115.130 161.245 115.455 161.705 ;
        RECT 115.975 161.075 116.255 161.535 ;
        RECT 115.130 160.855 116.255 161.075 ;
        RECT 114.575 159.895 114.855 160.565 ;
        RECT 115.130 160.395 115.580 160.855 ;
        RECT 116.445 160.685 116.845 161.535 ;
        RECT 117.245 161.245 117.515 161.705 ;
        RECT 117.685 161.075 117.970 161.535 ;
        RECT 115.025 160.065 115.580 160.395 ;
        RECT 115.750 160.125 116.845 160.685 ;
        RECT 115.130 159.955 115.580 160.065 ;
        RECT 114.575 159.325 114.960 159.895 ;
        RECT 115.130 159.785 116.255 159.955 ;
        RECT 115.130 159.155 115.455 159.615 ;
        RECT 115.975 159.325 116.255 159.785 ;
        RECT 116.445 159.325 116.845 160.125 ;
        RECT 117.015 160.855 117.970 161.075 ;
        RECT 117.015 159.955 117.225 160.855 ;
        RECT 117.395 160.125 118.085 160.685 ;
        RECT 118.255 160.615 119.465 161.705 ;
        RECT 118.255 160.075 118.775 160.615 ;
        RECT 117.015 159.785 117.970 159.955 ;
        RECT 118.945 159.905 119.465 160.445 ;
        RECT 117.245 159.155 117.515 159.615 ;
        RECT 117.685 159.325 117.970 159.785 ;
        RECT 118.255 159.155 119.465 159.905 ;
        RECT 71.250 158.985 119.550 159.155 ;
        RECT 71.335 158.235 72.545 158.985 ;
        RECT 72.715 158.440 78.060 158.985 ;
        RECT 71.335 157.695 71.855 158.235 ;
        RECT 72.025 157.525 72.545 158.065 ;
        RECT 74.300 157.610 74.640 158.440 ;
        RECT 78.235 158.215 80.825 158.985 ;
        RECT 81.505 158.595 81.835 158.985 ;
        RECT 82.005 158.415 82.175 158.735 ;
        RECT 82.345 158.595 82.675 158.985 ;
        RECT 83.090 158.585 84.045 158.755 ;
        RECT 81.455 158.245 83.705 158.415 ;
        RECT 71.335 156.435 72.545 157.525 ;
        RECT 76.120 156.870 76.470 158.120 ;
        RECT 78.235 157.695 79.445 158.215 ;
        RECT 79.615 157.525 80.825 158.045 ;
        RECT 72.715 156.435 78.060 156.870 ;
        RECT 78.235 156.435 80.825 157.525 ;
        RECT 81.455 157.285 81.625 158.245 ;
        RECT 81.795 157.625 82.040 158.075 ;
        RECT 82.210 157.795 82.760 157.995 ;
        RECT 82.930 157.825 83.305 157.995 ;
        RECT 82.930 157.625 83.100 157.825 ;
        RECT 83.475 157.745 83.705 158.245 ;
        RECT 81.795 157.455 83.100 157.625 ;
        RECT 83.875 157.705 84.045 158.585 ;
        RECT 84.215 158.150 84.505 158.985 ;
        RECT 84.675 158.150 84.965 158.985 ;
        RECT 85.135 158.585 86.090 158.755 ;
        RECT 86.505 158.595 86.835 158.985 ;
        RECT 85.135 157.705 85.305 158.585 ;
        RECT 87.005 158.415 87.175 158.735 ;
        RECT 87.345 158.595 87.675 158.985 ;
        RECT 87.945 158.595 88.275 158.985 ;
        RECT 88.445 158.415 88.615 158.735 ;
        RECT 88.785 158.595 89.115 158.985 ;
        RECT 89.530 158.585 90.485 158.755 ;
        RECT 85.475 158.245 87.725 158.415 ;
        RECT 85.475 157.745 85.705 158.245 ;
        RECT 85.875 157.825 86.250 157.995 ;
        RECT 83.875 157.535 84.505 157.705 ;
        RECT 81.455 156.605 81.835 157.285 ;
        RECT 82.425 156.435 82.595 157.285 ;
        RECT 82.765 157.115 84.005 157.285 ;
        RECT 82.765 156.605 83.095 157.115 ;
        RECT 83.265 156.435 83.435 156.945 ;
        RECT 83.605 156.605 84.005 157.115 ;
        RECT 84.185 156.605 84.505 157.535 ;
        RECT 84.675 157.535 85.305 157.705 ;
        RECT 86.080 157.625 86.250 157.825 ;
        RECT 86.420 157.795 86.970 157.995 ;
        RECT 87.140 157.625 87.385 158.075 ;
        RECT 84.675 156.605 84.995 157.535 ;
        RECT 86.080 157.455 87.385 157.625 ;
        RECT 87.555 157.285 87.725 158.245 ;
        RECT 85.175 157.115 86.415 157.285 ;
        RECT 85.175 156.605 85.575 157.115 ;
        RECT 85.745 156.435 85.915 156.945 ;
        RECT 86.085 156.605 86.415 157.115 ;
        RECT 86.585 156.435 86.755 157.285 ;
        RECT 87.345 156.605 87.725 157.285 ;
        RECT 87.895 158.245 90.145 158.415 ;
        RECT 87.895 157.285 88.065 158.245 ;
        RECT 88.235 157.625 88.480 158.075 ;
        RECT 88.650 157.795 89.200 157.995 ;
        RECT 89.370 157.825 89.745 157.995 ;
        RECT 89.370 157.625 89.540 157.825 ;
        RECT 89.915 157.745 90.145 158.245 ;
        RECT 88.235 157.455 89.540 157.625 ;
        RECT 90.315 157.705 90.485 158.585 ;
        RECT 90.655 158.150 90.945 158.985 ;
        RECT 91.690 158.355 91.975 158.815 ;
        RECT 92.145 158.525 92.415 158.985 ;
        RECT 91.690 158.185 92.645 158.355 ;
        RECT 90.315 157.535 90.945 157.705 ;
        RECT 87.895 156.605 88.275 157.285 ;
        RECT 88.865 156.435 89.035 157.285 ;
        RECT 89.205 157.115 90.445 157.285 ;
        RECT 89.205 156.605 89.535 157.115 ;
        RECT 89.705 156.435 89.875 156.945 ;
        RECT 90.045 156.605 90.445 157.115 ;
        RECT 90.625 156.605 90.945 157.535 ;
        RECT 91.575 157.455 92.265 158.015 ;
        RECT 92.435 157.285 92.645 158.185 ;
        RECT 91.690 157.065 92.645 157.285 ;
        RECT 92.815 158.015 93.215 158.815 ;
        RECT 93.405 158.355 93.685 158.815 ;
        RECT 94.205 158.525 94.530 158.985 ;
        RECT 93.405 158.185 94.530 158.355 ;
        RECT 94.700 158.245 95.085 158.815 ;
        RECT 94.080 158.075 94.530 158.185 ;
        RECT 92.815 157.455 93.910 158.015 ;
        RECT 94.080 157.745 94.635 158.075 ;
        RECT 91.690 156.605 91.975 157.065 ;
        RECT 92.145 156.435 92.415 156.895 ;
        RECT 92.815 156.605 93.215 157.455 ;
        RECT 94.080 157.285 94.530 157.745 ;
        RECT 94.805 157.575 95.085 158.245 ;
        RECT 95.255 158.215 96.925 158.985 ;
        RECT 97.095 158.260 97.385 158.985 ;
        RECT 97.555 158.215 101.065 158.985 ;
        RECT 95.255 157.695 96.005 158.215 ;
        RECT 93.405 157.065 94.530 157.285 ;
        RECT 93.405 156.605 93.685 157.065 ;
        RECT 94.205 156.435 94.530 156.895 ;
        RECT 94.700 156.605 95.085 157.575 ;
        RECT 96.175 157.525 96.925 158.045 ;
        RECT 97.555 157.695 99.205 158.215 ;
        RECT 101.695 158.185 102.035 158.815 ;
        RECT 102.325 158.525 102.495 158.985 ;
        RECT 102.765 158.355 103.095 158.800 ;
        RECT 95.255 156.435 96.925 157.525 ;
        RECT 97.095 156.435 97.385 157.600 ;
        RECT 99.375 157.525 101.065 158.045 ;
        RECT 97.555 156.435 101.065 157.525 ;
        RECT 101.695 157.615 101.965 158.185 ;
        RECT 102.345 158.165 103.095 158.355 ;
        RECT 103.265 158.335 103.435 158.655 ;
        RECT 103.660 158.525 103.990 158.985 ;
        RECT 104.190 158.335 104.520 158.815 ;
        RECT 104.735 158.525 105.065 158.985 ;
        RECT 105.235 158.335 105.565 158.815 ;
        RECT 103.265 158.165 105.565 158.335 ;
        RECT 102.345 157.995 102.715 158.165 ;
        RECT 102.135 157.785 102.715 157.995 ;
        RECT 102.885 157.785 103.305 157.995 ;
        RECT 102.455 157.615 102.715 157.785 ;
        RECT 101.695 156.605 102.220 157.615 ;
        RECT 102.455 157.325 103.205 157.615 ;
        RECT 102.455 156.435 102.785 157.155 ;
        RECT 102.955 156.605 103.205 157.325 ;
        RECT 103.475 156.680 103.805 157.995 ;
        RECT 104.015 156.680 104.345 157.995 ;
        RECT 104.515 156.680 104.885 157.995 ;
        RECT 105.095 157.745 105.605 157.995 ;
        RECT 105.215 156.435 105.545 157.555 ;
        RECT 106.295 156.605 106.555 158.815 ;
        RECT 106.805 158.525 106.975 158.985 ;
        RECT 107.145 158.645 108.140 158.815 ;
        RECT 108.670 158.655 108.840 158.815 ;
        RECT 107.145 158.355 107.315 158.645 ;
        RECT 107.970 158.485 108.140 158.645 ;
        RECT 108.310 158.485 108.840 158.655 ;
        RECT 106.745 158.185 107.315 158.355 ;
        RECT 107.485 158.305 107.660 158.475 ;
        RECT 106.745 157.405 106.915 158.185 ;
        RECT 107.485 158.145 107.900 158.305 ;
        RECT 107.490 158.135 107.900 158.145 ;
        RECT 107.225 157.795 107.680 157.965 ;
        RECT 106.745 157.235 107.395 157.405 ;
        RECT 108.310 157.315 108.480 158.485 ;
        RECT 109.185 158.415 109.360 158.745 ;
        RECT 109.530 158.605 109.860 158.985 ;
        RECT 108.650 158.135 108.890 158.305 ;
        RECT 106.725 156.435 107.055 156.815 ;
        RECT 107.225 156.775 107.395 157.235 ;
        RECT 107.695 157.085 108.480 157.315 ;
        RECT 107.695 156.945 108.025 157.085 ;
        RECT 108.720 156.935 108.890 158.135 ;
        RECT 109.185 157.965 109.355 158.415 ;
        RECT 110.130 158.355 110.375 158.775 ;
        RECT 110.550 158.525 110.720 158.985 ;
        RECT 110.890 158.645 112.490 158.815 ;
        RECT 110.890 158.605 111.245 158.645 ;
        RECT 111.480 158.355 111.650 158.475 ;
        RECT 110.130 158.185 111.650 158.355 ;
        RECT 111.480 158.145 111.650 158.185 ;
        RECT 111.820 158.225 112.150 158.475 ;
        RECT 112.320 158.275 112.490 158.645 ;
        RECT 112.780 158.265 113.070 158.985 ;
        RECT 113.780 158.645 114.855 158.815 ;
        RECT 111.820 158.150 112.135 158.225 ;
        RECT 109.065 157.795 109.355 157.965 ;
        RECT 108.180 156.775 108.510 156.815 ;
        RECT 107.225 156.605 108.510 156.775 ;
        RECT 108.680 156.605 108.890 156.935 ;
        RECT 109.185 156.935 109.355 157.795 ;
        RECT 109.525 157.395 109.815 158.075 ;
        RECT 110.290 157.625 110.620 158.015 ;
        RECT 110.265 157.455 110.620 157.625 ;
        RECT 110.290 157.395 110.620 157.455 ;
        RECT 110.825 157.625 111.070 158.015 ;
        RECT 111.465 157.965 111.795 157.975 ;
        RECT 111.410 157.805 111.795 157.965 ;
        RECT 111.410 157.795 111.580 157.805 ;
        RECT 111.965 157.625 112.135 158.150 ;
        RECT 110.825 157.455 111.125 157.625 ;
        RECT 111.375 157.455 112.135 157.625 ;
        RECT 110.825 157.395 111.070 157.455 ;
        RECT 110.140 156.985 111.205 157.155 ;
        RECT 109.185 156.605 109.370 156.935 ;
        RECT 109.540 156.435 109.890 156.815 ;
        RECT 110.140 156.605 110.310 156.985 ;
        RECT 110.480 156.435 110.810 156.815 ;
        RECT 111.035 156.775 111.205 156.985 ;
        RECT 111.375 156.945 111.705 157.455 ;
        RECT 111.875 156.775 112.045 157.285 ;
        RECT 112.305 157.075 112.605 158.075 ;
        RECT 113.250 157.965 113.610 158.640 ;
        RECT 113.780 158.310 113.950 158.645 ;
        RECT 114.120 158.305 114.460 158.475 ;
        RECT 114.170 158.135 114.460 158.305 ;
        RECT 114.685 158.435 114.855 158.645 ;
        RECT 115.025 158.605 115.355 158.985 ;
        RECT 115.525 158.435 115.695 158.810 ;
        RECT 114.685 158.265 115.695 158.435 ;
        RECT 113.250 157.785 113.790 157.965 ;
        RECT 113.250 157.675 113.610 157.785 ;
        RECT 112.805 157.445 113.610 157.675 ;
        RECT 114.290 157.615 114.460 158.135 ;
        RECT 115.955 158.215 117.625 158.985 ;
        RECT 118.255 158.235 119.465 158.985 ;
        RECT 113.825 157.445 114.460 157.615 ;
        RECT 114.630 157.455 115.065 158.075 ;
        RECT 115.375 157.625 115.720 158.075 ;
        RECT 115.955 157.695 116.705 158.215 ;
        RECT 115.375 157.455 115.725 157.625 ;
        RECT 116.875 157.525 117.625 158.045 ;
        RECT 111.035 156.605 112.045 156.775 ;
        RECT 112.305 156.435 112.635 156.815 ;
        RECT 112.805 156.605 113.155 157.445 ;
        RECT 113.325 156.775 113.495 157.275 ;
        RECT 113.825 157.115 113.995 157.445 ;
        RECT 113.665 156.945 113.995 157.115 ;
        RECT 114.165 157.105 115.695 157.275 ;
        RECT 114.165 156.945 114.335 157.105 ;
        RECT 114.685 156.775 114.855 156.935 ;
        RECT 113.325 156.605 114.855 156.775 ;
        RECT 115.025 156.435 115.355 156.815 ;
        RECT 115.525 156.605 115.695 157.105 ;
        RECT 115.955 156.435 117.625 157.525 ;
        RECT 118.255 157.525 118.775 158.065 ;
        RECT 118.945 157.695 119.465 158.235 ;
        RECT 118.255 156.435 119.465 157.525 ;
        RECT 71.250 156.265 119.550 156.435 ;
        RECT 71.335 155.175 72.545 156.265 ;
        RECT 73.640 155.595 73.895 156.095 ;
        RECT 74.065 155.765 74.395 156.265 ;
        RECT 73.640 155.425 74.390 155.595 ;
        RECT 71.335 154.465 71.855 155.005 ;
        RECT 72.025 154.635 72.545 155.175 ;
        RECT 73.640 154.605 73.990 155.255 ;
        RECT 71.335 153.715 72.545 154.465 ;
        RECT 74.160 154.435 74.390 155.425 ;
        RECT 73.640 154.265 74.390 154.435 ;
        RECT 73.640 153.975 73.895 154.265 ;
        RECT 74.065 153.715 74.395 154.095 ;
        RECT 74.565 153.975 74.735 156.095 ;
        RECT 74.905 155.295 75.230 156.080 ;
        RECT 75.400 155.805 75.650 156.265 ;
        RECT 75.820 155.765 76.070 156.095 ;
        RECT 76.285 155.765 76.965 156.095 ;
        RECT 75.820 155.635 75.990 155.765 ;
        RECT 75.595 155.465 75.990 155.635 ;
        RECT 74.965 154.245 75.425 155.295 ;
        RECT 75.595 154.105 75.765 155.465 ;
        RECT 76.160 155.205 76.625 155.595 ;
        RECT 75.935 154.395 76.285 155.015 ;
        RECT 76.455 154.615 76.625 155.205 ;
        RECT 76.795 154.985 76.965 155.765 ;
        RECT 77.135 155.665 77.305 156.005 ;
        RECT 77.540 155.835 77.870 156.265 ;
        RECT 78.040 155.665 78.210 156.005 ;
        RECT 78.505 155.805 78.875 156.265 ;
        RECT 77.135 155.495 78.210 155.665 ;
        RECT 79.045 155.635 79.215 156.095 ;
        RECT 79.450 155.755 80.320 156.095 ;
        RECT 80.490 155.805 80.740 156.265 ;
        RECT 78.655 155.465 79.215 155.635 ;
        RECT 78.655 155.325 78.825 155.465 ;
        RECT 77.325 155.155 78.825 155.325 ;
        RECT 79.520 155.295 79.980 155.585 ;
        RECT 76.795 154.815 78.485 154.985 ;
        RECT 76.455 154.395 76.810 154.615 ;
        RECT 76.980 154.105 77.150 154.815 ;
        RECT 77.355 154.395 78.145 154.645 ;
        RECT 78.315 154.635 78.485 154.815 ;
        RECT 78.655 154.465 78.825 155.155 ;
        RECT 75.095 153.715 75.425 154.075 ;
        RECT 75.595 153.935 76.090 154.105 ;
        RECT 76.295 153.935 77.150 154.105 ;
        RECT 78.025 153.715 78.355 154.175 ;
        RECT 78.565 154.075 78.825 154.465 ;
        RECT 79.015 155.285 79.980 155.295 ;
        RECT 80.150 155.375 80.320 155.755 ;
        RECT 80.910 155.715 81.080 156.005 ;
        RECT 81.260 155.885 81.590 156.265 ;
        RECT 80.910 155.545 81.710 155.715 ;
        RECT 79.015 155.125 79.690 155.285 ;
        RECT 80.150 155.205 81.370 155.375 ;
        RECT 79.015 154.335 79.225 155.125 ;
        RECT 80.150 155.115 80.320 155.205 ;
        RECT 79.395 154.335 79.745 154.955 ;
        RECT 79.915 154.945 80.320 155.115 ;
        RECT 79.915 154.165 80.085 154.945 ;
        RECT 80.255 154.495 80.475 154.775 ;
        RECT 80.655 154.665 81.195 155.035 ;
        RECT 81.540 154.955 81.710 155.545 ;
        RECT 81.930 155.125 82.235 156.265 ;
        RECT 82.405 155.075 82.660 155.955 ;
        RECT 82.835 155.175 84.045 156.265 ;
        RECT 81.540 154.925 82.280 154.955 ;
        RECT 80.255 154.325 80.785 154.495 ;
        RECT 78.565 153.905 78.915 154.075 ;
        RECT 79.135 153.885 80.085 154.165 ;
        RECT 80.255 153.715 80.445 154.155 ;
        RECT 80.615 154.095 80.785 154.325 ;
        RECT 80.955 154.265 81.195 154.665 ;
        RECT 81.365 154.625 82.280 154.925 ;
        RECT 81.365 154.450 81.690 154.625 ;
        RECT 81.365 154.095 81.685 154.450 ;
        RECT 82.450 154.425 82.660 155.075 ;
        RECT 80.615 153.925 81.685 154.095 ;
        RECT 81.930 153.715 82.235 154.175 ;
        RECT 82.405 153.895 82.660 154.425 ;
        RECT 82.835 154.465 83.355 155.005 ;
        RECT 83.525 154.635 84.045 155.175 ;
        RECT 84.215 155.100 84.505 156.265 ;
        RECT 84.675 155.125 85.060 156.095 ;
        RECT 85.230 155.805 85.555 156.265 ;
        RECT 86.075 155.635 86.355 156.095 ;
        RECT 85.230 155.415 86.355 155.635 ;
        RECT 82.835 153.715 84.045 154.465 ;
        RECT 84.675 154.455 84.955 155.125 ;
        RECT 85.230 154.955 85.680 155.415 ;
        RECT 86.545 155.245 86.945 156.095 ;
        RECT 87.345 155.805 87.615 156.265 ;
        RECT 87.785 155.635 88.070 156.095 ;
        RECT 85.125 154.625 85.680 154.955 ;
        RECT 85.850 154.685 86.945 155.245 ;
        RECT 85.230 154.515 85.680 154.625 ;
        RECT 84.215 153.715 84.505 154.440 ;
        RECT 84.675 153.885 85.060 154.455 ;
        RECT 85.230 154.345 86.355 154.515 ;
        RECT 85.230 153.715 85.555 154.175 ;
        RECT 86.075 153.885 86.355 154.345 ;
        RECT 86.545 153.885 86.945 154.685 ;
        RECT 87.115 155.415 88.070 155.635 ;
        RECT 87.115 154.515 87.325 155.415 ;
        RECT 87.495 154.685 88.185 155.245 ;
        RECT 88.355 155.125 88.740 156.095 ;
        RECT 88.910 155.805 89.235 156.265 ;
        RECT 89.755 155.635 90.035 156.095 ;
        RECT 88.910 155.415 90.035 155.635 ;
        RECT 87.115 154.345 88.070 154.515 ;
        RECT 87.345 153.715 87.615 154.175 ;
        RECT 87.785 153.885 88.070 154.345 ;
        RECT 88.355 154.455 88.635 155.125 ;
        RECT 88.910 154.955 89.360 155.415 ;
        RECT 90.225 155.245 90.625 156.095 ;
        RECT 91.025 155.805 91.295 156.265 ;
        RECT 91.465 155.635 91.750 156.095 ;
        RECT 88.805 154.625 89.360 154.955 ;
        RECT 89.530 154.685 90.625 155.245 ;
        RECT 88.910 154.515 89.360 154.625 ;
        RECT 88.355 153.885 88.740 154.455 ;
        RECT 88.910 154.345 90.035 154.515 ;
        RECT 88.910 153.715 89.235 154.175 ;
        RECT 89.755 153.885 90.035 154.345 ;
        RECT 90.225 153.885 90.625 154.685 ;
        RECT 90.795 155.415 91.750 155.635 ;
        RECT 92.040 155.595 92.295 156.095 ;
        RECT 92.465 155.765 92.795 156.265 ;
        RECT 92.040 155.425 92.790 155.595 ;
        RECT 90.795 154.515 91.005 155.415 ;
        RECT 91.175 154.685 91.865 155.245 ;
        RECT 92.040 154.605 92.390 155.255 ;
        RECT 90.795 154.345 91.750 154.515 ;
        RECT 92.560 154.435 92.790 155.425 ;
        RECT 91.025 153.715 91.295 154.175 ;
        RECT 91.465 153.885 91.750 154.345 ;
        RECT 92.040 154.265 92.790 154.435 ;
        RECT 92.040 153.975 92.295 154.265 ;
        RECT 92.465 153.715 92.795 154.095 ;
        RECT 92.965 153.975 93.135 156.095 ;
        RECT 93.305 155.295 93.630 156.080 ;
        RECT 93.800 155.805 94.050 156.265 ;
        RECT 94.220 155.765 94.470 156.095 ;
        RECT 94.685 155.765 95.365 156.095 ;
        RECT 94.220 155.635 94.390 155.765 ;
        RECT 93.995 155.465 94.390 155.635 ;
        RECT 93.365 154.245 93.825 155.295 ;
        RECT 93.995 154.105 94.165 155.465 ;
        RECT 94.560 155.205 95.025 155.595 ;
        RECT 94.335 154.395 94.685 155.015 ;
        RECT 94.855 154.615 95.025 155.205 ;
        RECT 95.195 154.985 95.365 155.765 ;
        RECT 95.535 155.665 95.705 156.005 ;
        RECT 95.940 155.835 96.270 156.265 ;
        RECT 96.440 155.665 96.610 156.005 ;
        RECT 96.905 155.805 97.275 156.265 ;
        RECT 95.535 155.495 96.610 155.665 ;
        RECT 97.445 155.635 97.615 156.095 ;
        RECT 97.850 155.755 98.720 156.095 ;
        RECT 98.890 155.805 99.140 156.265 ;
        RECT 97.055 155.465 97.615 155.635 ;
        RECT 97.055 155.325 97.225 155.465 ;
        RECT 95.725 155.155 97.225 155.325 ;
        RECT 97.920 155.295 98.380 155.585 ;
        RECT 95.195 154.815 96.885 154.985 ;
        RECT 94.855 154.395 95.210 154.615 ;
        RECT 95.380 154.105 95.550 154.815 ;
        RECT 95.755 154.395 96.545 154.645 ;
        RECT 96.715 154.635 96.885 154.815 ;
        RECT 97.055 154.465 97.225 155.155 ;
        RECT 93.495 153.715 93.825 154.075 ;
        RECT 93.995 153.935 94.490 154.105 ;
        RECT 94.695 153.935 95.550 154.105 ;
        RECT 96.425 153.715 96.755 154.175 ;
        RECT 96.965 154.075 97.225 154.465 ;
        RECT 97.415 155.285 98.380 155.295 ;
        RECT 98.550 155.375 98.720 155.755 ;
        RECT 99.310 155.715 99.480 156.005 ;
        RECT 99.660 155.885 99.990 156.265 ;
        RECT 99.310 155.545 100.110 155.715 ;
        RECT 97.415 155.125 98.090 155.285 ;
        RECT 98.550 155.205 99.770 155.375 ;
        RECT 97.415 154.335 97.625 155.125 ;
        RECT 98.550 155.115 98.720 155.205 ;
        RECT 97.795 154.335 98.145 154.955 ;
        RECT 98.315 154.945 98.720 155.115 ;
        RECT 98.315 154.165 98.485 154.945 ;
        RECT 98.655 154.495 98.875 154.775 ;
        RECT 99.055 154.665 99.595 155.035 ;
        RECT 99.940 154.955 100.110 155.545 ;
        RECT 100.330 155.125 100.635 156.265 ;
        RECT 100.805 155.075 101.060 155.955 ;
        RECT 101.325 155.595 101.495 156.095 ;
        RECT 101.665 155.765 101.995 156.265 ;
        RECT 101.325 155.425 101.990 155.595 ;
        RECT 99.940 154.925 100.680 154.955 ;
        RECT 98.655 154.325 99.185 154.495 ;
        RECT 96.965 153.905 97.315 154.075 ;
        RECT 97.535 153.885 98.485 154.165 ;
        RECT 98.655 153.715 98.845 154.155 ;
        RECT 99.015 154.095 99.185 154.325 ;
        RECT 99.355 154.265 99.595 154.665 ;
        RECT 99.765 154.625 100.680 154.925 ;
        RECT 99.765 154.450 100.090 154.625 ;
        RECT 99.765 154.095 100.085 154.450 ;
        RECT 100.850 154.425 101.060 155.075 ;
        RECT 101.240 154.605 101.590 155.255 ;
        RECT 101.760 154.435 101.990 155.425 ;
        RECT 99.015 153.925 100.085 154.095 ;
        RECT 100.330 153.715 100.635 154.175 ;
        RECT 100.805 153.895 101.060 154.425 ;
        RECT 101.325 154.265 101.990 154.435 ;
        RECT 101.325 153.975 101.495 154.265 ;
        RECT 101.665 153.715 101.995 154.095 ;
        RECT 102.165 153.975 102.350 156.095 ;
        RECT 102.590 155.805 102.855 156.265 ;
        RECT 103.025 155.670 103.275 156.095 ;
        RECT 103.485 155.820 104.590 155.990 ;
        RECT 102.970 155.540 103.275 155.670 ;
        RECT 102.520 154.345 102.800 155.295 ;
        RECT 102.970 154.435 103.140 155.540 ;
        RECT 103.310 154.755 103.550 155.350 ;
        RECT 103.720 155.285 104.250 155.650 ;
        RECT 103.720 154.585 103.890 155.285 ;
        RECT 104.420 155.205 104.590 155.820 ;
        RECT 104.760 155.465 104.930 156.265 ;
        RECT 105.100 155.765 105.350 156.095 ;
        RECT 105.575 155.795 106.460 155.965 ;
        RECT 104.420 155.115 104.930 155.205 ;
        RECT 102.970 154.305 103.195 154.435 ;
        RECT 103.365 154.365 103.890 154.585 ;
        RECT 104.060 154.945 104.930 155.115 ;
        RECT 102.605 153.715 102.855 154.175 ;
        RECT 103.025 154.165 103.195 154.305 ;
        RECT 104.060 154.165 104.230 154.945 ;
        RECT 104.760 154.875 104.930 154.945 ;
        RECT 104.440 154.695 104.640 154.725 ;
        RECT 105.100 154.695 105.270 155.765 ;
        RECT 105.440 154.875 105.630 155.595 ;
        RECT 104.440 154.395 105.270 154.695 ;
        RECT 105.800 154.665 106.120 155.625 ;
        RECT 103.025 153.995 103.360 154.165 ;
        RECT 103.555 153.995 104.230 154.165 ;
        RECT 104.550 153.715 104.920 154.215 ;
        RECT 105.100 154.165 105.270 154.395 ;
        RECT 105.655 154.335 106.120 154.665 ;
        RECT 106.290 154.955 106.460 155.795 ;
        RECT 106.640 155.765 106.955 156.265 ;
        RECT 107.185 155.535 107.525 156.095 ;
        RECT 106.630 155.160 107.525 155.535 ;
        RECT 107.695 155.255 107.865 156.265 ;
        RECT 107.335 154.955 107.525 155.160 ;
        RECT 108.035 155.205 108.365 156.050 ;
        RECT 108.035 155.125 108.425 155.205 ;
        RECT 108.655 155.125 108.865 156.265 ;
        RECT 108.210 155.075 108.425 155.125 ;
        RECT 106.290 154.625 107.165 154.955 ;
        RECT 107.335 154.625 108.085 154.955 ;
        RECT 106.290 154.165 106.460 154.625 ;
        RECT 107.335 154.455 107.535 154.625 ;
        RECT 108.255 154.495 108.425 155.075 ;
        RECT 109.035 155.115 109.365 156.095 ;
        RECT 109.535 155.125 109.765 156.265 ;
        RECT 108.200 154.455 108.425 154.495 ;
        RECT 105.100 153.995 105.505 154.165 ;
        RECT 105.675 153.995 106.460 154.165 ;
        RECT 106.735 153.715 106.945 154.245 ;
        RECT 107.205 153.930 107.535 154.455 ;
        RECT 108.045 154.370 108.425 154.455 ;
        RECT 107.705 153.715 107.875 154.325 ;
        RECT 108.045 153.935 108.375 154.370 ;
        RECT 108.655 153.715 108.865 154.535 ;
        RECT 109.035 154.515 109.285 155.115 ;
        RECT 109.975 155.100 110.265 156.265 ;
        RECT 110.985 155.595 111.155 156.095 ;
        RECT 111.325 155.765 111.655 156.265 ;
        RECT 110.985 155.425 111.650 155.595 ;
        RECT 109.455 154.705 109.785 154.955 ;
        RECT 110.900 154.605 111.250 155.255 ;
        RECT 109.035 153.885 109.365 154.515 ;
        RECT 109.535 153.715 109.765 154.535 ;
        RECT 109.975 153.715 110.265 154.440 ;
        RECT 111.420 154.435 111.650 155.425 ;
        RECT 110.985 154.265 111.650 154.435 ;
        RECT 110.985 153.975 111.155 154.265 ;
        RECT 111.325 153.715 111.655 154.095 ;
        RECT 111.825 153.975 112.010 156.095 ;
        RECT 112.250 155.805 112.515 156.265 ;
        RECT 112.685 155.670 112.935 156.095 ;
        RECT 113.145 155.820 114.250 155.990 ;
        RECT 112.630 155.540 112.935 155.670 ;
        RECT 112.180 154.345 112.460 155.295 ;
        RECT 112.630 154.435 112.800 155.540 ;
        RECT 112.970 154.755 113.210 155.350 ;
        RECT 113.380 155.285 113.910 155.650 ;
        RECT 113.380 154.585 113.550 155.285 ;
        RECT 114.080 155.205 114.250 155.820 ;
        RECT 114.420 155.465 114.590 156.265 ;
        RECT 114.760 155.765 115.010 156.095 ;
        RECT 115.235 155.795 116.120 155.965 ;
        RECT 114.080 155.115 114.590 155.205 ;
        RECT 112.630 154.305 112.855 154.435 ;
        RECT 113.025 154.365 113.550 154.585 ;
        RECT 113.720 154.945 114.590 155.115 ;
        RECT 112.265 153.715 112.515 154.175 ;
        RECT 112.685 154.165 112.855 154.305 ;
        RECT 113.720 154.165 113.890 154.945 ;
        RECT 114.420 154.875 114.590 154.945 ;
        RECT 114.100 154.695 114.300 154.725 ;
        RECT 114.760 154.695 114.930 155.765 ;
        RECT 115.100 154.875 115.290 155.595 ;
        RECT 114.100 154.395 114.930 154.695 ;
        RECT 115.460 154.665 115.780 155.625 ;
        RECT 112.685 153.995 113.020 154.165 ;
        RECT 113.215 153.995 113.890 154.165 ;
        RECT 114.210 153.715 114.580 154.215 ;
        RECT 114.760 154.165 114.930 154.395 ;
        RECT 115.315 154.335 115.780 154.665 ;
        RECT 115.950 154.955 116.120 155.795 ;
        RECT 116.300 155.765 116.615 156.265 ;
        RECT 116.845 155.535 117.185 156.095 ;
        RECT 116.290 155.160 117.185 155.535 ;
        RECT 117.355 155.255 117.525 156.265 ;
        RECT 116.995 154.955 117.185 155.160 ;
        RECT 117.695 155.205 118.025 156.050 ;
        RECT 117.695 155.125 118.085 155.205 ;
        RECT 117.870 155.075 118.085 155.125 ;
        RECT 115.950 154.625 116.825 154.955 ;
        RECT 116.995 154.625 117.745 154.955 ;
        RECT 115.950 154.165 116.120 154.625 ;
        RECT 116.995 154.455 117.195 154.625 ;
        RECT 117.915 154.495 118.085 155.075 ;
        RECT 118.255 155.175 119.465 156.265 ;
        RECT 118.255 154.635 118.775 155.175 ;
        RECT 117.860 154.455 118.085 154.495 ;
        RECT 118.945 154.465 119.465 155.005 ;
        RECT 114.760 153.995 115.165 154.165 ;
        RECT 115.335 153.995 116.120 154.165 ;
        RECT 116.395 153.715 116.605 154.245 ;
        RECT 116.865 153.930 117.195 154.455 ;
        RECT 117.705 154.370 118.085 154.455 ;
        RECT 117.365 153.715 117.535 154.325 ;
        RECT 117.705 153.935 118.035 154.370 ;
        RECT 118.255 153.715 119.465 154.465 ;
        RECT 71.250 153.545 119.550 153.715 ;
        RECT 17.610 152.920 17.985 153.265 ;
        RECT 20.630 152.940 20.965 153.285 ;
        RECT 71.335 152.795 72.545 153.545 ;
        RECT 18.300 152.355 21.080 152.525 ;
        RECT 18.300 151.885 18.470 152.355 ;
        RECT 18.090 151.375 18.590 151.885 ;
        RECT 14.840 148.000 16.515 148.550 ;
        RECT 18.300 148.000 18.470 151.375 ;
        RECT 18.960 151.145 19.130 152.185 ;
        RECT 19.400 151.145 19.570 152.355 ;
        RECT 19.840 151.145 20.010 152.185 ;
        RECT 20.470 151.145 20.640 152.185 ;
        RECT 20.910 151.145 21.080 152.355 ;
        RECT 71.335 152.255 71.855 152.795 ;
        RECT 72.715 152.775 76.225 153.545 ;
        RECT 76.395 152.795 77.605 153.545 ;
        RECT 77.775 152.805 78.160 153.375 ;
        RECT 78.330 153.085 78.655 153.545 ;
        RECT 79.175 152.915 79.455 153.375 ;
        RECT 21.350 151.145 21.520 152.185 ;
        RECT 72.025 152.085 72.545 152.625 ;
        RECT 72.715 152.255 74.365 152.775 ;
        RECT 74.535 152.085 76.225 152.605 ;
        RECT 76.395 152.255 76.915 152.795 ;
        RECT 77.085 152.085 77.605 152.625 ;
        RECT 71.335 150.995 72.545 152.085 ;
        RECT 72.715 150.995 76.225 152.085 ;
        RECT 76.395 150.995 77.605 152.085 ;
        RECT 77.775 152.135 78.055 152.805 ;
        RECT 78.330 152.745 79.455 152.915 ;
        RECT 78.330 152.635 78.780 152.745 ;
        RECT 78.225 152.305 78.780 152.635 ;
        RECT 79.645 152.575 80.045 153.375 ;
        RECT 80.445 153.085 80.715 153.545 ;
        RECT 80.885 152.915 81.170 153.375 ;
        RECT 77.775 151.165 78.160 152.135 ;
        RECT 78.330 151.845 78.780 152.305 ;
        RECT 78.950 152.015 80.045 152.575 ;
        RECT 78.330 151.625 79.455 151.845 ;
        RECT 78.330 150.995 78.655 151.455 ;
        RECT 79.175 151.165 79.455 151.625 ;
        RECT 79.645 151.165 80.045 152.015 ;
        RECT 80.215 152.745 81.170 152.915 ;
        RECT 80.215 151.845 80.425 152.745 ;
        RECT 81.455 152.710 81.745 153.545 ;
        RECT 81.915 153.145 82.870 153.315 ;
        RECT 83.285 153.155 83.615 153.545 ;
        RECT 80.595 152.015 81.285 152.575 ;
        RECT 81.915 152.265 82.085 153.145 ;
        RECT 83.785 152.975 83.955 153.295 ;
        RECT 84.125 153.155 84.455 153.545 ;
        RECT 82.255 152.805 84.505 152.975 ;
        RECT 82.255 152.305 82.485 152.805 ;
        RECT 82.655 152.385 83.030 152.555 ;
        RECT 81.455 152.095 82.085 152.265 ;
        RECT 82.860 152.185 83.030 152.385 ;
        RECT 83.200 152.355 83.750 152.555 ;
        RECT 83.920 152.185 84.165 152.635 ;
        RECT 80.215 151.625 81.170 151.845 ;
        RECT 80.445 150.995 80.715 151.455 ;
        RECT 80.885 151.165 81.170 151.625 ;
        RECT 81.455 151.165 81.775 152.095 ;
        RECT 82.860 152.015 84.165 152.185 ;
        RECT 84.335 151.845 84.505 152.805 ;
        RECT 84.675 152.775 87.265 153.545 ;
        RECT 87.985 153.065 88.285 153.545 ;
        RECT 88.455 152.895 88.715 153.350 ;
        RECT 88.885 153.065 89.145 153.545 ;
        RECT 89.325 152.895 89.585 153.350 ;
        RECT 89.755 153.065 90.005 153.545 ;
        RECT 90.185 152.895 90.445 153.350 ;
        RECT 90.615 153.065 90.865 153.545 ;
        RECT 91.045 152.895 91.305 153.350 ;
        RECT 91.475 153.065 91.720 153.545 ;
        RECT 91.890 152.895 92.165 153.350 ;
        RECT 92.335 153.065 92.580 153.545 ;
        RECT 92.750 152.895 93.010 153.350 ;
        RECT 93.180 153.065 93.440 153.545 ;
        RECT 93.610 152.895 93.870 153.350 ;
        RECT 94.040 153.065 94.300 153.545 ;
        RECT 94.470 152.895 94.730 153.350 ;
        RECT 94.900 152.985 95.160 153.545 ;
        RECT 84.675 152.255 85.885 152.775 ;
        RECT 87.985 152.725 94.730 152.895 ;
        RECT 86.055 152.085 87.265 152.605 ;
        RECT 81.955 151.675 83.195 151.845 ;
        RECT 81.955 151.165 82.355 151.675 ;
        RECT 82.525 150.995 82.695 151.505 ;
        RECT 82.865 151.165 83.195 151.675 ;
        RECT 83.365 150.995 83.535 151.845 ;
        RECT 84.125 151.165 84.505 151.845 ;
        RECT 84.675 150.995 87.265 152.085 ;
        RECT 87.985 152.135 89.150 152.725 ;
        RECT 95.330 152.555 95.580 153.365 ;
        RECT 95.760 153.020 96.020 153.545 ;
        RECT 96.190 152.555 96.440 153.365 ;
        RECT 96.620 153.035 96.925 153.545 ;
        RECT 89.320 152.305 96.440 152.555 ;
        RECT 96.610 152.305 96.925 152.865 ;
        RECT 97.095 152.820 97.385 153.545 ;
        RECT 97.555 152.775 100.145 153.545 ;
        RECT 100.775 152.805 101.265 153.375 ;
        RECT 101.435 152.975 101.665 153.375 ;
        RECT 101.835 153.145 102.255 153.545 ;
        RECT 102.425 152.975 102.595 153.375 ;
        RECT 101.435 152.805 102.595 152.975 ;
        RECT 102.765 152.805 103.215 153.545 ;
        RECT 103.385 152.805 103.825 153.365 ;
        RECT 104.085 152.995 104.255 153.285 ;
        RECT 104.425 153.165 104.755 153.545 ;
        RECT 104.085 152.825 104.750 152.995 ;
        RECT 87.985 151.910 94.730 152.135 ;
        RECT 87.985 150.995 88.255 151.740 ;
        RECT 88.425 151.170 88.715 151.910 ;
        RECT 89.325 151.895 94.730 151.910 ;
        RECT 88.885 151.000 89.140 151.725 ;
        RECT 89.325 151.170 89.585 151.895 ;
        RECT 89.755 151.000 90.000 151.725 ;
        RECT 90.185 151.170 90.445 151.895 ;
        RECT 90.615 151.000 90.860 151.725 ;
        RECT 91.045 151.170 91.305 151.895 ;
        RECT 91.475 151.000 91.720 151.725 ;
        RECT 91.890 151.170 92.150 151.895 ;
        RECT 92.320 151.000 92.580 151.725 ;
        RECT 92.750 151.170 93.010 151.895 ;
        RECT 93.180 151.000 93.440 151.725 ;
        RECT 93.610 151.170 93.870 151.895 ;
        RECT 94.040 151.000 94.300 151.725 ;
        RECT 94.470 151.170 94.730 151.895 ;
        RECT 94.900 151.000 95.160 151.795 ;
        RECT 95.330 151.170 95.580 152.305 ;
        RECT 88.885 150.995 95.160 151.000 ;
        RECT 95.760 150.995 96.020 151.805 ;
        RECT 96.195 151.165 96.440 152.305 ;
        RECT 97.555 152.255 98.765 152.775 ;
        RECT 96.620 150.995 96.915 151.805 ;
        RECT 97.095 150.995 97.385 152.160 ;
        RECT 98.935 152.085 100.145 152.605 ;
        RECT 97.555 150.995 100.145 152.085 ;
        RECT 100.775 152.135 100.945 152.805 ;
        RECT 101.115 152.305 101.520 152.635 ;
        RECT 100.775 151.965 101.545 152.135 ;
        RECT 100.785 150.995 101.115 151.795 ;
        RECT 101.295 151.335 101.545 151.965 ;
        RECT 101.735 151.505 101.985 152.635 ;
        RECT 102.185 152.305 102.430 152.635 ;
        RECT 102.615 152.355 103.005 152.635 ;
        RECT 102.185 151.505 102.385 152.305 ;
        RECT 103.175 152.185 103.345 152.635 ;
        RECT 102.555 152.015 103.345 152.185 ;
        RECT 102.555 151.335 102.725 152.015 ;
        RECT 101.295 151.165 102.725 151.335 ;
        RECT 102.895 150.995 103.210 151.845 ;
        RECT 103.515 151.795 103.825 152.805 ;
        RECT 104.000 152.005 104.350 152.655 ;
        RECT 104.520 151.835 104.750 152.825 ;
        RECT 103.385 151.165 103.825 151.795 ;
        RECT 104.085 151.665 104.750 151.835 ;
        RECT 104.085 151.165 104.255 151.665 ;
        RECT 104.425 150.995 104.755 151.495 ;
        RECT 104.925 151.165 105.110 153.285 ;
        RECT 105.365 153.085 105.615 153.545 ;
        RECT 105.785 153.095 106.120 153.265 ;
        RECT 106.315 153.095 106.990 153.265 ;
        RECT 105.785 152.955 105.955 153.095 ;
        RECT 105.280 151.965 105.560 152.915 ;
        RECT 105.730 152.825 105.955 152.955 ;
        RECT 105.730 151.720 105.900 152.825 ;
        RECT 106.125 152.675 106.650 152.895 ;
        RECT 106.070 151.910 106.310 152.505 ;
        RECT 106.480 151.975 106.650 152.675 ;
        RECT 106.820 152.315 106.990 153.095 ;
        RECT 107.310 153.045 107.680 153.545 ;
        RECT 107.860 153.095 108.265 153.265 ;
        RECT 108.435 153.095 109.220 153.265 ;
        RECT 107.860 152.865 108.030 153.095 ;
        RECT 107.200 152.565 108.030 152.865 ;
        RECT 108.415 152.595 108.880 152.925 ;
        RECT 107.200 152.535 107.400 152.565 ;
        RECT 107.520 152.315 107.690 152.385 ;
        RECT 106.820 152.145 107.690 152.315 ;
        RECT 107.180 152.055 107.690 152.145 ;
        RECT 105.730 151.590 106.035 151.720 ;
        RECT 106.480 151.610 107.010 151.975 ;
        RECT 105.350 150.995 105.615 151.455 ;
        RECT 105.785 151.165 106.035 151.590 ;
        RECT 107.180 151.440 107.350 152.055 ;
        RECT 106.245 151.270 107.350 151.440 ;
        RECT 107.520 150.995 107.690 151.795 ;
        RECT 107.860 151.495 108.030 152.565 ;
        RECT 108.200 151.665 108.390 152.385 ;
        RECT 108.560 151.635 108.880 152.595 ;
        RECT 109.050 152.635 109.220 153.095 ;
        RECT 109.495 153.015 109.705 153.545 ;
        RECT 109.965 152.805 110.295 153.330 ;
        RECT 110.465 152.935 110.635 153.545 ;
        RECT 110.805 152.890 111.135 153.325 ;
        RECT 111.930 152.915 112.215 153.375 ;
        RECT 112.385 153.085 112.655 153.545 ;
        RECT 110.805 152.805 111.185 152.890 ;
        RECT 110.095 152.635 110.295 152.805 ;
        RECT 110.960 152.765 111.185 152.805 ;
        RECT 109.050 152.305 109.925 152.635 ;
        RECT 110.095 152.305 110.845 152.635 ;
        RECT 107.860 151.165 108.110 151.495 ;
        RECT 109.050 151.465 109.220 152.305 ;
        RECT 110.095 152.100 110.285 152.305 ;
        RECT 111.015 152.185 111.185 152.765 ;
        RECT 111.930 152.745 112.885 152.915 ;
        RECT 110.970 152.135 111.185 152.185 ;
        RECT 109.390 151.725 110.285 152.100 ;
        RECT 110.795 152.055 111.185 152.135 ;
        RECT 108.335 151.295 109.220 151.465 ;
        RECT 109.400 150.995 109.715 151.495 ;
        RECT 109.945 151.165 110.285 151.725 ;
        RECT 110.455 150.995 110.625 152.005 ;
        RECT 110.795 151.210 111.125 152.055 ;
        RECT 111.815 152.015 112.505 152.575 ;
        RECT 112.675 151.845 112.885 152.745 ;
        RECT 111.930 151.625 112.885 151.845 ;
        RECT 113.055 152.575 113.455 153.375 ;
        RECT 113.645 152.915 113.925 153.375 ;
        RECT 114.445 153.085 114.770 153.545 ;
        RECT 113.645 152.745 114.770 152.915 ;
        RECT 114.940 152.805 115.325 153.375 ;
        RECT 114.320 152.635 114.770 152.745 ;
        RECT 113.055 152.015 114.150 152.575 ;
        RECT 114.320 152.305 114.875 152.635 ;
        RECT 111.930 151.165 112.215 151.625 ;
        RECT 112.385 150.995 112.655 151.455 ;
        RECT 113.055 151.165 113.455 152.015 ;
        RECT 114.320 151.845 114.770 152.305 ;
        RECT 115.045 152.135 115.325 152.805 ;
        RECT 115.495 152.795 116.705 153.545 ;
        RECT 116.875 152.870 117.135 153.375 ;
        RECT 117.315 153.165 117.645 153.545 ;
        RECT 117.825 152.995 117.995 153.375 ;
        RECT 115.495 152.255 116.015 152.795 ;
        RECT 113.645 151.625 114.770 151.845 ;
        RECT 113.645 151.165 113.925 151.625 ;
        RECT 114.445 150.995 114.770 151.455 ;
        RECT 114.940 151.165 115.325 152.135 ;
        RECT 116.185 152.085 116.705 152.625 ;
        RECT 115.495 150.995 116.705 152.085 ;
        RECT 116.875 152.070 117.055 152.870 ;
        RECT 117.330 152.825 117.995 152.995 ;
        RECT 117.330 152.570 117.500 152.825 ;
        RECT 118.255 152.795 119.465 153.545 ;
        RECT 117.225 152.240 117.500 152.570 ;
        RECT 117.725 152.275 118.065 152.645 ;
        RECT 117.330 152.095 117.500 152.240 ;
        RECT 116.875 151.165 117.145 152.070 ;
        RECT 117.330 151.925 118.005 152.095 ;
        RECT 117.315 150.995 117.645 151.755 ;
        RECT 117.825 151.165 118.005 151.925 ;
        RECT 118.255 152.085 118.775 152.625 ;
        RECT 118.945 152.255 119.465 152.795 ;
        RECT 118.255 150.995 119.465 152.085 ;
        RECT 71.250 150.825 119.550 150.995 ;
        RECT 21.130 150.240 21.300 150.570 ;
        RECT 71.335 149.735 72.545 150.825 ;
        RECT 72.715 150.390 78.060 150.825 ;
        RECT 71.335 149.025 71.855 149.565 ;
        RECT 72.025 149.195 72.545 149.735 ;
        RECT 71.335 148.275 72.545 149.025 ;
        RECT 74.300 148.820 74.640 149.650 ;
        RECT 76.120 149.140 76.470 150.390 ;
        RECT 78.235 149.735 80.825 150.825 ;
        RECT 78.235 149.045 79.445 149.565 ;
        RECT 79.615 149.215 80.825 149.735 ;
        RECT 80.995 149.750 81.265 150.655 ;
        RECT 81.435 150.065 81.765 150.825 ;
        RECT 81.945 149.895 82.115 150.655 ;
        RECT 72.715 148.275 78.060 148.820 ;
        RECT 78.235 148.275 80.825 149.045 ;
        RECT 80.995 148.950 81.165 149.750 ;
        RECT 81.450 149.725 82.115 149.895 ;
        RECT 82.375 149.735 84.045 150.825 ;
        RECT 81.450 149.580 81.620 149.725 ;
        RECT 81.335 149.250 81.620 149.580 ;
        RECT 81.450 148.995 81.620 149.250 ;
        RECT 81.855 149.175 82.185 149.545 ;
        RECT 82.375 149.045 83.125 149.565 ;
        RECT 83.295 149.215 84.045 149.735 ;
        RECT 84.215 149.660 84.505 150.825 ;
        RECT 84.680 150.155 84.935 150.655 ;
        RECT 85.105 150.325 85.435 150.825 ;
        RECT 84.680 149.985 85.430 150.155 ;
        RECT 84.680 149.165 85.030 149.815 ;
        RECT 80.995 148.445 81.255 148.950 ;
        RECT 81.450 148.825 82.115 148.995 ;
        RECT 81.435 148.275 81.765 148.655 ;
        RECT 81.945 148.445 82.115 148.825 ;
        RECT 82.375 148.275 84.045 149.045 ;
        RECT 84.215 148.275 84.505 149.000 ;
        RECT 85.200 148.995 85.430 149.985 ;
        RECT 84.680 148.825 85.430 148.995 ;
        RECT 84.680 148.535 84.935 148.825 ;
        RECT 85.105 148.275 85.435 148.655 ;
        RECT 85.605 148.535 85.775 150.655 ;
        RECT 85.945 149.855 86.270 150.640 ;
        RECT 86.440 150.365 86.690 150.825 ;
        RECT 86.860 150.325 87.110 150.655 ;
        RECT 87.325 150.325 88.005 150.655 ;
        RECT 86.860 150.195 87.030 150.325 ;
        RECT 86.635 150.025 87.030 150.195 ;
        RECT 86.005 148.805 86.465 149.855 ;
        RECT 86.635 148.665 86.805 150.025 ;
        RECT 87.200 149.765 87.665 150.155 ;
        RECT 86.975 148.955 87.325 149.575 ;
        RECT 87.495 149.175 87.665 149.765 ;
        RECT 87.835 149.545 88.005 150.325 ;
        RECT 88.175 150.225 88.345 150.565 ;
        RECT 88.580 150.395 88.910 150.825 ;
        RECT 89.080 150.225 89.250 150.565 ;
        RECT 89.545 150.365 89.915 150.825 ;
        RECT 88.175 150.055 89.250 150.225 ;
        RECT 90.085 150.195 90.255 150.655 ;
        RECT 90.490 150.315 91.360 150.655 ;
        RECT 91.530 150.365 91.780 150.825 ;
        RECT 89.695 150.025 90.255 150.195 ;
        RECT 89.695 149.885 89.865 150.025 ;
        RECT 88.365 149.715 89.865 149.885 ;
        RECT 90.560 149.855 91.020 150.145 ;
        RECT 87.835 149.375 89.525 149.545 ;
        RECT 87.495 148.955 87.850 149.175 ;
        RECT 88.020 148.665 88.190 149.375 ;
        RECT 88.395 148.955 89.185 149.205 ;
        RECT 89.355 149.195 89.525 149.375 ;
        RECT 89.695 149.025 89.865 149.715 ;
        RECT 86.135 148.275 86.465 148.635 ;
        RECT 86.635 148.495 87.130 148.665 ;
        RECT 87.335 148.495 88.190 148.665 ;
        RECT 89.065 148.275 89.395 148.735 ;
        RECT 89.605 148.635 89.865 149.025 ;
        RECT 90.055 149.845 91.020 149.855 ;
        RECT 91.190 149.935 91.360 150.315 ;
        RECT 91.950 150.275 92.120 150.565 ;
        RECT 92.300 150.445 92.630 150.825 ;
        RECT 91.950 150.105 92.750 150.275 ;
        RECT 90.055 149.685 90.730 149.845 ;
        RECT 91.190 149.765 92.410 149.935 ;
        RECT 90.055 148.895 90.265 149.685 ;
        RECT 91.190 149.675 91.360 149.765 ;
        RECT 90.435 148.895 90.785 149.515 ;
        RECT 90.955 149.505 91.360 149.675 ;
        RECT 90.955 148.725 91.125 149.505 ;
        RECT 91.295 149.055 91.515 149.335 ;
        RECT 91.695 149.225 92.235 149.595 ;
        RECT 92.580 149.515 92.750 150.105 ;
        RECT 92.970 149.685 93.275 150.825 ;
        RECT 93.445 149.635 93.700 150.515 ;
        RECT 93.875 149.735 96.465 150.825 ;
        RECT 92.580 149.485 93.320 149.515 ;
        RECT 91.295 148.885 91.825 149.055 ;
        RECT 89.605 148.465 89.955 148.635 ;
        RECT 90.175 148.445 91.125 148.725 ;
        RECT 91.295 148.275 91.485 148.715 ;
        RECT 91.655 148.655 91.825 148.885 ;
        RECT 91.995 148.825 92.235 149.225 ;
        RECT 92.405 149.185 93.320 149.485 ;
        RECT 92.405 149.010 92.730 149.185 ;
        RECT 92.405 148.655 92.725 149.010 ;
        RECT 93.490 148.985 93.700 149.635 ;
        RECT 91.655 148.485 92.725 148.655 ;
        RECT 92.970 148.275 93.275 148.735 ;
        RECT 93.445 148.455 93.700 148.985 ;
        RECT 93.875 149.045 95.085 149.565 ;
        RECT 95.255 149.215 96.465 149.735 ;
        RECT 97.095 149.660 97.385 150.825 ;
        RECT 97.555 150.390 102.900 150.825 ;
        RECT 93.875 148.275 96.465 149.045 ;
        RECT 97.095 148.275 97.385 149.000 ;
        RECT 99.140 148.820 99.480 149.650 ;
        RECT 100.960 149.140 101.310 150.390 ;
        RECT 103.075 149.735 104.285 150.825 ;
        RECT 103.075 149.025 103.595 149.565 ;
        RECT 103.765 149.195 104.285 149.735 ;
        RECT 104.545 149.895 104.715 150.655 ;
        RECT 104.895 150.065 105.225 150.825 ;
        RECT 104.545 149.725 105.210 149.895 ;
        RECT 105.395 149.750 105.665 150.655 ;
        RECT 105.040 149.580 105.210 149.725 ;
        RECT 104.475 149.175 104.805 149.545 ;
        RECT 105.040 149.250 105.325 149.580 ;
        RECT 97.555 148.275 102.900 148.820 ;
        RECT 103.075 148.275 104.285 149.025 ;
        RECT 105.040 148.995 105.210 149.250 ;
        RECT 104.545 148.825 105.210 148.995 ;
        RECT 105.495 148.950 105.665 149.750 ;
        RECT 104.545 148.445 104.715 148.825 ;
        RECT 104.895 148.275 105.225 148.655 ;
        RECT 105.405 148.445 105.665 148.950 ;
        RECT 105.835 150.025 106.275 150.655 ;
        RECT 105.835 149.015 106.145 150.025 ;
        RECT 106.450 149.975 106.765 150.825 ;
        RECT 106.935 150.485 108.365 150.655 ;
        RECT 106.935 149.805 107.105 150.485 ;
        RECT 106.315 149.635 107.105 149.805 ;
        RECT 106.315 149.185 106.485 149.635 ;
        RECT 107.275 149.515 107.475 150.315 ;
        RECT 106.655 149.185 107.045 149.465 ;
        RECT 107.230 149.185 107.475 149.515 ;
        RECT 107.675 149.185 107.925 150.315 ;
        RECT 108.115 149.855 108.365 150.485 ;
        RECT 108.545 150.025 108.875 150.825 ;
        RECT 108.115 149.685 108.885 149.855 ;
        RECT 108.140 149.185 108.545 149.515 ;
        RECT 108.715 149.015 108.885 149.685 ;
        RECT 109.975 149.660 110.265 150.825 ;
        RECT 110.435 149.685 110.820 150.655 ;
        RECT 110.990 150.365 111.315 150.825 ;
        RECT 111.835 150.195 112.115 150.655 ;
        RECT 110.990 149.975 112.115 150.195 ;
        RECT 105.835 148.455 106.275 149.015 ;
        RECT 106.445 148.275 106.895 149.015 ;
        RECT 107.065 148.845 108.225 149.015 ;
        RECT 107.065 148.445 107.235 148.845 ;
        RECT 107.405 148.275 107.825 148.675 ;
        RECT 107.995 148.445 108.225 148.845 ;
        RECT 108.395 148.445 108.885 149.015 ;
        RECT 110.435 149.015 110.715 149.685 ;
        RECT 110.990 149.515 111.440 149.975 ;
        RECT 112.305 149.805 112.705 150.655 ;
        RECT 113.105 150.365 113.375 150.825 ;
        RECT 113.545 150.195 113.830 150.655 ;
        RECT 110.885 149.185 111.440 149.515 ;
        RECT 111.610 149.245 112.705 149.805 ;
        RECT 110.990 149.075 111.440 149.185 ;
        RECT 109.975 148.275 110.265 149.000 ;
        RECT 110.435 148.445 110.820 149.015 ;
        RECT 110.990 148.905 112.115 149.075 ;
        RECT 110.990 148.275 111.315 148.735 ;
        RECT 111.835 148.445 112.115 148.905 ;
        RECT 112.305 148.445 112.705 149.245 ;
        RECT 112.875 149.975 113.830 150.195 ;
        RECT 112.875 149.075 113.085 149.975 ;
        RECT 113.255 149.245 113.945 149.805 ;
        RECT 114.575 149.685 114.960 150.655 ;
        RECT 115.130 150.365 115.455 150.825 ;
        RECT 115.975 150.195 116.255 150.655 ;
        RECT 115.130 149.975 116.255 150.195 ;
        RECT 112.875 148.905 113.830 149.075 ;
        RECT 113.105 148.275 113.375 148.735 ;
        RECT 113.545 148.445 113.830 148.905 ;
        RECT 114.575 149.015 114.855 149.685 ;
        RECT 115.130 149.515 115.580 149.975 ;
        RECT 116.445 149.805 116.845 150.655 ;
        RECT 117.245 150.365 117.515 150.825 ;
        RECT 117.685 150.195 117.970 150.655 ;
        RECT 115.025 149.185 115.580 149.515 ;
        RECT 115.750 149.245 116.845 149.805 ;
        RECT 115.130 149.075 115.580 149.185 ;
        RECT 114.575 148.445 114.960 149.015 ;
        RECT 115.130 148.905 116.255 149.075 ;
        RECT 115.130 148.275 115.455 148.735 ;
        RECT 115.975 148.445 116.255 148.905 ;
        RECT 116.445 148.445 116.845 149.245 ;
        RECT 117.015 149.975 117.970 150.195 ;
        RECT 117.015 149.075 117.225 149.975 ;
        RECT 117.395 149.245 118.085 149.805 ;
        RECT 118.255 149.735 119.465 150.825 ;
        RECT 118.255 149.195 118.775 149.735 ;
        RECT 117.015 148.905 117.970 149.075 ;
        RECT 118.945 149.025 119.465 149.565 ;
        RECT 117.245 148.275 117.515 148.735 ;
        RECT 117.685 148.445 117.970 148.905 ;
        RECT 118.255 148.275 119.465 149.025 ;
        RECT 71.250 148.105 119.550 148.275 ;
        RECT 14.840 147.830 18.470 148.000 ;
        RECT 14.840 147.275 16.515 147.830 ;
        RECT 18.300 139.270 18.470 147.830 ;
        RECT 13.095 139.100 18.470 139.270 ;
        RECT 13.095 137.140 13.265 139.100 ;
        RECT 14.535 137.510 30.905 137.680 ;
        RECT 12.885 136.820 13.270 137.140 ;
        RECT 11.850 136.010 12.280 136.080 ;
        RECT 12.655 136.010 12.825 136.540 ;
        RECT 11.850 135.835 12.825 136.010 ;
        RECT 11.850 135.700 12.280 135.835 ;
        RECT 12.655 135.500 12.825 135.835 ;
        RECT 13.095 135.500 13.265 136.820 ;
        RECT 12.570 132.520 12.920 134.680 ;
        RECT 14.535 132.230 14.705 137.510 ;
        RECT 17.210 136.155 17.380 136.665 ;
        RECT 17.210 135.985 18.960 136.155 ;
        RECT 17.210 133.585 17.380 135.985 ;
        RECT 17.920 135.475 18.250 135.645 ;
        RECT 17.780 134.265 17.950 135.305 ;
        RECT 18.220 134.955 18.390 135.305 ;
        RECT 18.790 134.955 18.960 135.985 ;
        RECT 19.240 135.985 20.990 136.155 ;
        RECT 19.240 134.955 19.410 135.985 ;
        RECT 19.950 135.475 20.280 135.645 ;
        RECT 19.810 134.955 19.980 135.305 ;
        RECT 18.190 134.675 19.980 134.955 ;
        RECT 18.220 134.265 18.390 134.675 ;
        RECT 17.920 133.925 18.250 134.095 ;
        RECT 18.790 133.585 18.960 134.675 ;
        RECT 19.240 133.585 19.410 134.675 ;
        RECT 19.810 134.265 19.980 134.675 ;
        RECT 20.250 134.265 20.420 135.305 ;
        RECT 19.950 133.925 20.280 134.095 ;
        RECT 20.820 133.585 20.990 135.985 ;
        RECT 21.270 135.985 23.020 136.155 ;
        RECT 21.270 133.585 21.440 135.985 ;
        RECT 21.980 135.475 22.310 135.645 ;
        RECT 21.840 134.265 22.010 135.305 ;
        RECT 22.280 134.265 22.450 135.305 ;
        RECT 21.980 133.925 22.310 134.095 ;
        RECT 22.850 133.595 23.020 135.985 ;
        RECT 23.300 135.995 25.050 136.165 ;
        RECT 23.300 133.595 23.470 135.995 ;
        RECT 24.010 135.485 24.340 135.655 ;
        RECT 23.870 134.275 24.040 135.315 ;
        RECT 24.310 134.275 24.480 135.315 ;
        RECT 24.010 133.935 24.340 134.105 ;
        RECT 24.880 133.595 25.050 135.995 ;
        RECT 25.320 135.995 27.070 136.165 ;
        RECT 25.320 133.595 25.490 135.995 ;
        RECT 26.030 135.485 26.360 135.655 ;
        RECT 25.890 134.275 26.060 135.315 ;
        RECT 26.330 134.935 26.500 135.315 ;
        RECT 26.900 134.935 27.070 135.995 ;
        RECT 27.345 135.990 29.095 136.160 ;
        RECT 27.345 134.935 27.515 135.990 ;
        RECT 28.055 135.480 28.385 135.650 ;
        RECT 27.915 134.935 28.085 135.310 ;
        RECT 26.310 134.655 28.100 134.935 ;
        RECT 26.330 134.275 26.500 134.655 ;
        RECT 26.030 133.935 26.360 134.105 ;
        RECT 26.900 133.595 27.070 134.655 ;
        RECT 27.345 133.595 27.515 134.655 ;
        RECT 27.915 134.270 28.085 134.655 ;
        RECT 28.355 134.270 28.525 135.310 ;
        RECT 28.055 133.930 28.385 134.100 ;
        RECT 22.850 133.590 27.515 133.595 ;
        RECT 28.925 133.590 29.095 135.990 ;
        RECT 22.850 133.585 29.095 133.590 ;
        RECT 17.210 133.425 29.095 133.585 ;
        RECT 17.210 133.415 23.020 133.425 ;
        RECT 27.345 133.420 29.095 133.425 ;
        RECT 30.735 132.230 30.905 137.510 ;
        RECT 14.535 132.060 30.905 132.230 ;
        RECT 12.570 129.860 12.920 132.020 ;
        RECT 17.390 114.950 17.765 115.295 ;
        RECT 20.410 114.970 20.745 115.315 ;
        RECT 18.080 114.385 20.860 114.555 ;
        RECT 18.080 113.915 18.250 114.385 ;
        RECT 17.870 113.405 18.370 113.915 ;
        RECT 14.230 109.455 15.745 109.985 ;
        RECT 18.080 109.455 18.250 113.405 ;
        RECT 18.740 113.175 18.910 114.215 ;
        RECT 19.180 113.175 19.350 114.385 ;
        RECT 19.620 113.175 19.790 114.215 ;
        RECT 20.250 113.175 20.420 114.215 ;
        RECT 20.690 113.175 20.860 114.385 ;
        RECT 21.130 113.175 21.300 114.215 ;
        RECT 20.910 112.270 21.080 112.600 ;
        RECT 14.230 109.285 18.250 109.455 ;
        RECT 14.230 108.720 15.745 109.285 ;
        RECT 18.080 101.300 18.250 109.285 ;
        RECT 12.875 101.130 18.250 101.300 ;
        RECT 12.875 99.170 13.045 101.130 ;
        RECT 14.315 99.540 30.685 99.710 ;
        RECT 12.665 98.850 13.050 99.170 ;
        RECT 11.630 98.040 12.060 98.110 ;
        RECT 12.435 98.040 12.605 98.570 ;
        RECT 11.630 97.865 12.605 98.040 ;
        RECT 11.630 97.730 12.060 97.865 ;
        RECT 12.435 97.530 12.605 97.865 ;
        RECT 12.875 97.530 13.045 98.850 ;
        RECT 12.350 94.550 12.700 96.710 ;
        RECT 14.315 94.260 14.485 99.540 ;
        RECT 16.990 98.185 17.160 98.695 ;
        RECT 16.990 98.015 18.740 98.185 ;
        RECT 16.990 95.615 17.160 98.015 ;
        RECT 17.700 97.505 18.030 97.675 ;
        RECT 17.560 96.295 17.730 97.335 ;
        RECT 18.000 96.985 18.170 97.335 ;
        RECT 18.570 96.985 18.740 98.015 ;
        RECT 19.020 98.015 20.770 98.185 ;
        RECT 19.020 96.985 19.190 98.015 ;
        RECT 19.730 97.505 20.060 97.675 ;
        RECT 19.590 96.985 19.760 97.335 ;
        RECT 17.970 96.705 19.760 96.985 ;
        RECT 18.000 96.295 18.170 96.705 ;
        RECT 17.700 95.955 18.030 96.125 ;
        RECT 18.570 95.615 18.740 96.705 ;
        RECT 19.020 95.615 19.190 96.705 ;
        RECT 19.590 96.295 19.760 96.705 ;
        RECT 20.030 96.295 20.200 97.335 ;
        RECT 19.730 95.955 20.060 96.125 ;
        RECT 20.600 95.615 20.770 98.015 ;
        RECT 21.050 98.015 22.800 98.185 ;
        RECT 21.050 95.615 21.220 98.015 ;
        RECT 21.760 97.505 22.090 97.675 ;
        RECT 21.620 96.295 21.790 97.335 ;
        RECT 22.060 96.295 22.230 97.335 ;
        RECT 21.760 95.955 22.090 96.125 ;
        RECT 22.630 95.625 22.800 98.015 ;
        RECT 23.080 98.025 24.830 98.195 ;
        RECT 23.080 95.625 23.250 98.025 ;
        RECT 23.790 97.515 24.120 97.685 ;
        RECT 23.650 96.305 23.820 97.345 ;
        RECT 24.090 96.305 24.260 97.345 ;
        RECT 23.790 95.965 24.120 96.135 ;
        RECT 24.660 95.625 24.830 98.025 ;
        RECT 25.100 98.025 26.850 98.195 ;
        RECT 25.100 95.625 25.270 98.025 ;
        RECT 25.810 97.515 26.140 97.685 ;
        RECT 25.670 96.305 25.840 97.345 ;
        RECT 26.110 96.965 26.280 97.345 ;
        RECT 26.680 96.965 26.850 98.025 ;
        RECT 27.125 98.020 28.875 98.190 ;
        RECT 27.125 96.965 27.295 98.020 ;
        RECT 27.835 97.510 28.165 97.680 ;
        RECT 27.695 96.965 27.865 97.340 ;
        RECT 26.090 96.685 27.880 96.965 ;
        RECT 26.110 96.305 26.280 96.685 ;
        RECT 25.810 95.965 26.140 96.135 ;
        RECT 26.680 95.625 26.850 96.685 ;
        RECT 27.125 95.625 27.295 96.685 ;
        RECT 27.695 96.300 27.865 96.685 ;
        RECT 28.135 96.300 28.305 97.340 ;
        RECT 27.835 95.960 28.165 96.130 ;
        RECT 22.630 95.620 27.295 95.625 ;
        RECT 28.705 95.620 28.875 98.020 ;
        RECT 22.630 95.615 28.875 95.620 ;
        RECT 16.990 95.455 28.875 95.615 ;
        RECT 16.990 95.445 22.800 95.455 ;
        RECT 27.125 95.450 28.875 95.455 ;
        RECT 30.515 94.260 30.685 99.540 ;
        RECT 14.315 94.090 30.685 94.260 ;
        RECT 12.350 91.890 12.700 94.050 ;
        RECT 91.060 88.855 152.240 89.025 ;
        RECT 91.145 88.105 92.355 88.855 ;
        RECT 92.525 88.310 97.870 88.855 ;
        RECT 98.045 88.310 103.390 88.855 ;
        RECT 91.145 87.565 91.665 88.105 ;
        RECT 91.835 87.395 92.355 87.935 ;
        RECT 94.110 87.480 94.450 88.310 ;
        RECT 91.145 86.305 92.355 87.395 ;
        RECT 95.930 86.740 96.280 87.990 ;
        RECT 99.630 87.480 99.970 88.310 ;
        RECT 104.025 88.130 104.315 88.855 ;
        RECT 104.545 88.375 104.825 88.855 ;
        RECT 104.995 88.205 105.255 88.595 ;
        RECT 105.430 88.375 105.685 88.855 ;
        RECT 105.855 88.205 106.150 88.595 ;
        RECT 106.330 88.375 106.605 88.855 ;
        RECT 106.775 88.355 107.075 88.685 ;
        RECT 104.500 88.035 106.150 88.205 ;
        RECT 101.450 86.740 101.800 87.990 ;
        RECT 104.500 87.525 104.905 88.035 ;
        RECT 105.075 87.695 106.215 87.865 ;
        RECT 92.525 86.305 97.870 86.740 ;
        RECT 98.045 86.305 103.390 86.740 ;
        RECT 104.025 86.305 104.315 87.470 ;
        RECT 104.500 87.355 105.255 87.525 ;
        RECT 104.540 86.305 104.825 87.175 ;
        RECT 104.995 87.105 105.255 87.355 ;
        RECT 106.045 87.445 106.215 87.695 ;
        RECT 106.385 87.615 106.735 88.185 ;
        RECT 106.905 87.445 107.075 88.355 ;
        RECT 107.245 88.310 112.590 88.855 ;
        RECT 108.830 87.480 109.170 88.310 ;
        RECT 112.765 88.085 116.275 88.855 ;
        RECT 116.905 88.130 117.195 88.855 ;
        RECT 117.365 88.310 122.710 88.855 ;
        RECT 122.885 88.310 128.230 88.855 ;
        RECT 106.045 87.275 107.075 87.445 ;
        RECT 104.995 86.935 106.115 87.105 ;
        RECT 104.995 86.475 105.255 86.935 ;
        RECT 105.430 86.305 105.685 86.765 ;
        RECT 105.855 86.475 106.115 86.935 ;
        RECT 106.285 86.305 106.595 87.105 ;
        RECT 106.765 86.475 107.075 87.275 ;
        RECT 110.650 86.740 111.000 87.990 ;
        RECT 112.765 87.565 114.415 88.085 ;
        RECT 114.585 87.395 116.275 87.915 ;
        RECT 118.950 87.480 119.290 88.310 ;
        RECT 107.245 86.305 112.590 86.740 ;
        RECT 112.765 86.305 116.275 87.395 ;
        RECT 116.905 86.305 117.195 87.470 ;
        RECT 120.770 86.740 121.120 87.990 ;
        RECT 124.470 87.480 124.810 88.310 ;
        RECT 128.405 88.105 129.615 88.855 ;
        RECT 129.785 88.130 130.075 88.855 ;
        RECT 130.245 88.310 135.590 88.855 ;
        RECT 126.290 86.740 126.640 87.990 ;
        RECT 128.405 87.565 128.925 88.105 ;
        RECT 129.095 87.395 129.615 87.935 ;
        RECT 131.830 87.480 132.170 88.310 ;
        RECT 135.765 88.085 139.275 88.855 ;
        RECT 139.905 88.355 140.205 88.685 ;
        RECT 140.375 88.375 140.650 88.855 ;
        RECT 117.365 86.305 122.710 86.740 ;
        RECT 122.885 86.305 128.230 86.740 ;
        RECT 128.405 86.305 129.615 87.395 ;
        RECT 129.785 86.305 130.075 87.470 ;
        RECT 133.650 86.740 134.000 87.990 ;
        RECT 135.765 87.565 137.415 88.085 ;
        RECT 137.585 87.395 139.275 87.915 ;
        RECT 130.245 86.305 135.590 86.740 ;
        RECT 135.765 86.305 139.275 87.395 ;
        RECT 139.905 87.445 140.075 88.355 ;
        RECT 140.830 88.205 141.125 88.595 ;
        RECT 141.295 88.375 141.550 88.855 ;
        RECT 141.725 88.205 141.985 88.595 ;
        RECT 142.155 88.375 142.435 88.855 ;
        RECT 140.245 87.615 140.595 88.185 ;
        RECT 140.830 88.035 142.480 88.205 ;
        RECT 142.665 88.130 142.955 88.855 ;
        RECT 143.125 88.310 148.470 88.855 ;
        RECT 149.110 88.455 149.445 88.855 ;
        RECT 140.765 87.695 141.905 87.865 ;
        RECT 140.765 87.445 140.935 87.695 ;
        RECT 142.075 87.525 142.480 88.035 ;
        RECT 139.905 87.275 140.935 87.445 ;
        RECT 141.725 87.355 142.480 87.525 ;
        RECT 144.710 87.480 145.050 88.310 ;
        RECT 149.615 88.285 149.820 88.685 ;
        RECT 150.030 88.375 150.305 88.855 ;
        RECT 150.515 88.355 150.775 88.685 ;
        RECT 149.135 88.115 149.820 88.285 ;
        RECT 139.905 86.475 140.215 87.275 ;
        RECT 141.725 87.105 141.985 87.355 ;
        RECT 140.385 86.305 140.695 87.105 ;
        RECT 140.865 86.935 141.985 87.105 ;
        RECT 140.865 86.475 141.125 86.935 ;
        RECT 141.295 86.305 141.550 86.765 ;
        RECT 141.725 86.475 141.985 86.935 ;
        RECT 142.155 86.305 142.440 87.175 ;
        RECT 142.665 86.305 142.955 87.470 ;
        RECT 146.530 86.740 146.880 87.990 ;
        RECT 149.135 87.085 149.475 88.115 ;
        RECT 149.645 87.445 149.895 87.945 ;
        RECT 150.075 87.615 150.435 88.195 ;
        RECT 150.605 87.445 150.775 88.355 ;
        RECT 150.945 88.105 152.155 88.855 ;
        RECT 149.645 87.275 150.775 87.445 ;
        RECT 149.135 86.910 149.800 87.085 ;
        RECT 143.125 86.305 148.470 86.740 ;
        RECT 149.110 86.305 149.445 86.730 ;
        RECT 149.615 86.505 149.800 86.910 ;
        RECT 150.005 86.305 150.335 87.085 ;
        RECT 150.505 86.505 150.775 87.275 ;
        RECT 150.945 87.395 151.465 87.935 ;
        RECT 151.635 87.565 152.155 88.105 ;
        RECT 150.945 86.305 152.155 87.395 ;
        RECT 91.060 86.135 152.240 86.305 ;
        RECT 91.145 85.045 92.355 86.135 ;
        RECT 92.525 85.700 97.870 86.135 ;
        RECT 98.045 85.700 103.390 86.135 ;
        RECT 91.145 84.335 91.665 84.875 ;
        RECT 91.835 84.505 92.355 85.045 ;
        RECT 91.145 83.585 92.355 84.335 ;
        RECT 94.110 84.130 94.450 84.960 ;
        RECT 95.930 84.450 96.280 85.700 ;
        RECT 99.630 84.130 99.970 84.960 ;
        RECT 101.450 84.450 101.800 85.700 ;
        RECT 104.025 84.970 104.315 86.135 ;
        RECT 104.485 85.700 109.830 86.135 ;
        RECT 110.005 85.700 115.350 86.135 ;
        RECT 115.525 85.700 120.870 86.135 ;
        RECT 92.525 83.585 97.870 84.130 ;
        RECT 98.045 83.585 103.390 84.130 ;
        RECT 104.025 83.585 104.315 84.310 ;
        RECT 106.070 84.130 106.410 84.960 ;
        RECT 107.890 84.450 108.240 85.700 ;
        RECT 111.590 84.130 111.930 84.960 ;
        RECT 113.410 84.450 113.760 85.700 ;
        RECT 117.110 84.130 117.450 84.960 ;
        RECT 118.930 84.450 119.280 85.700 ;
        RECT 121.965 84.995 122.245 86.135 ;
        RECT 122.415 84.985 122.745 85.965 ;
        RECT 122.915 84.995 123.175 86.135 ;
        RECT 123.345 85.045 125.015 86.135 ;
        RECT 121.975 84.555 122.310 84.825 ;
        RECT 122.480 84.385 122.650 84.985 ;
        RECT 122.820 84.575 123.155 84.825 ;
        RECT 104.485 83.585 109.830 84.130 ;
        RECT 110.005 83.585 115.350 84.130 ;
        RECT 115.525 83.585 120.870 84.130 ;
        RECT 121.965 83.585 122.275 84.385 ;
        RECT 122.480 83.755 123.175 84.385 ;
        RECT 123.345 84.355 124.095 84.875 ;
        RECT 124.265 84.525 125.015 85.045 ;
        RECT 125.185 85.060 125.455 85.965 ;
        RECT 125.625 85.375 125.955 86.135 ;
        RECT 126.135 85.205 126.305 85.965 ;
        RECT 123.345 83.585 125.015 84.355 ;
        RECT 125.185 84.260 125.355 85.060 ;
        RECT 125.640 85.035 126.305 85.205 ;
        RECT 126.565 85.045 129.155 86.135 ;
        RECT 125.640 84.890 125.810 85.035 ;
        RECT 125.525 84.560 125.810 84.890 ;
        RECT 125.640 84.305 125.810 84.560 ;
        RECT 126.045 84.485 126.375 84.855 ;
        RECT 126.565 84.355 127.775 84.875 ;
        RECT 127.945 84.525 129.155 85.045 ;
        RECT 129.785 84.970 130.075 86.135 ;
        RECT 130.445 85.465 130.725 86.135 ;
        RECT 130.895 85.245 131.195 85.795 ;
        RECT 131.395 85.415 131.725 86.135 ;
        RECT 131.915 85.415 132.375 85.965 ;
        RECT 130.260 84.825 130.525 85.185 ;
        RECT 130.895 85.075 131.835 85.245 ;
        RECT 131.665 84.825 131.835 85.075 ;
        RECT 130.260 84.575 130.935 84.825 ;
        RECT 131.155 84.575 131.495 84.825 ;
        RECT 131.665 84.495 131.955 84.825 ;
        RECT 131.665 84.405 131.835 84.495 ;
        RECT 125.185 83.755 125.445 84.260 ;
        RECT 125.640 84.135 126.305 84.305 ;
        RECT 125.625 83.585 125.955 83.965 ;
        RECT 126.135 83.755 126.305 84.135 ;
        RECT 126.565 83.585 129.155 84.355 ;
        RECT 129.785 83.585 130.075 84.310 ;
        RECT 130.445 84.215 131.835 84.405 ;
        RECT 130.445 83.855 130.775 84.215 ;
        RECT 132.125 84.045 132.375 85.415 ;
        RECT 132.545 85.045 133.755 86.135 ;
        RECT 131.395 83.585 131.645 84.045 ;
        RECT 131.815 83.755 132.375 84.045 ;
        RECT 132.545 84.335 133.065 84.875 ;
        RECT 133.235 84.505 133.755 85.045 ;
        RECT 134.015 85.205 134.185 85.965 ;
        RECT 134.365 85.375 134.695 86.135 ;
        RECT 134.015 85.035 134.680 85.205 ;
        RECT 134.865 85.060 135.135 85.965 ;
        RECT 134.510 84.890 134.680 85.035 ;
        RECT 133.945 84.485 134.275 84.855 ;
        RECT 134.510 84.560 134.795 84.890 ;
        RECT 132.545 83.585 133.755 84.335 ;
        RECT 134.510 84.305 134.680 84.560 ;
        RECT 134.015 84.135 134.680 84.305 ;
        RECT 134.965 84.260 135.135 85.060 ;
        RECT 135.305 85.045 136.515 86.135 ;
        RECT 136.690 85.465 136.945 85.965 ;
        RECT 137.115 85.635 137.445 86.135 ;
        RECT 136.690 85.295 137.440 85.465 ;
        RECT 134.015 83.755 134.185 84.135 ;
        RECT 134.365 83.585 134.695 83.965 ;
        RECT 134.875 83.755 135.135 84.260 ;
        RECT 135.305 84.335 135.825 84.875 ;
        RECT 135.995 84.505 136.515 85.045 ;
        RECT 136.690 84.475 137.040 85.125 ;
        RECT 135.305 83.585 136.515 84.335 ;
        RECT 137.210 84.305 137.440 85.295 ;
        RECT 136.690 84.135 137.440 84.305 ;
        RECT 136.690 83.845 136.945 84.135 ;
        RECT 137.115 83.585 137.445 83.965 ;
        RECT 137.615 83.845 137.785 85.965 ;
        RECT 137.955 85.165 138.280 85.950 ;
        RECT 138.450 85.675 138.700 86.135 ;
        RECT 138.870 85.635 139.120 85.965 ;
        RECT 139.335 85.635 140.015 85.965 ;
        RECT 138.870 85.505 139.040 85.635 ;
        RECT 138.645 85.335 139.040 85.505 ;
        RECT 138.015 84.115 138.475 85.165 ;
        RECT 138.645 83.975 138.815 85.335 ;
        RECT 139.210 85.075 139.675 85.465 ;
        RECT 138.985 84.265 139.335 84.885 ;
        RECT 139.505 84.485 139.675 85.075 ;
        RECT 139.845 84.855 140.015 85.635 ;
        RECT 140.185 85.535 140.355 85.875 ;
        RECT 140.590 85.705 140.920 86.135 ;
        RECT 141.090 85.535 141.260 85.875 ;
        RECT 141.555 85.675 141.925 86.135 ;
        RECT 140.185 85.365 141.260 85.535 ;
        RECT 142.095 85.505 142.265 85.965 ;
        RECT 142.500 85.625 143.370 85.965 ;
        RECT 143.540 85.675 143.790 86.135 ;
        RECT 141.705 85.335 142.265 85.505 ;
        RECT 141.705 85.195 141.875 85.335 ;
        RECT 140.375 85.025 141.875 85.195 ;
        RECT 142.570 85.165 143.030 85.455 ;
        RECT 139.845 84.685 141.535 84.855 ;
        RECT 139.505 84.265 139.860 84.485 ;
        RECT 140.030 83.975 140.200 84.685 ;
        RECT 140.405 84.265 141.195 84.515 ;
        RECT 141.365 84.505 141.535 84.685 ;
        RECT 141.705 84.335 141.875 85.025 ;
        RECT 138.145 83.585 138.475 83.945 ;
        RECT 138.645 83.805 139.140 83.975 ;
        RECT 139.345 83.805 140.200 83.975 ;
        RECT 141.075 83.585 141.405 84.045 ;
        RECT 141.615 83.945 141.875 84.335 ;
        RECT 142.065 85.155 143.030 85.165 ;
        RECT 143.200 85.245 143.370 85.625 ;
        RECT 143.960 85.585 144.130 85.875 ;
        RECT 144.310 85.755 144.640 86.135 ;
        RECT 143.960 85.415 144.760 85.585 ;
        RECT 142.065 84.995 142.740 85.155 ;
        RECT 143.200 85.075 144.420 85.245 ;
        RECT 142.065 84.205 142.275 84.995 ;
        RECT 143.200 84.985 143.370 85.075 ;
        RECT 142.445 84.205 142.795 84.825 ;
        RECT 142.965 84.815 143.370 84.985 ;
        RECT 142.965 84.035 143.135 84.815 ;
        RECT 143.305 84.365 143.525 84.645 ;
        RECT 143.705 84.535 144.245 84.905 ;
        RECT 144.590 84.825 144.760 85.415 ;
        RECT 144.980 84.995 145.285 86.135 ;
        RECT 145.455 84.945 145.705 85.825 ;
        RECT 145.875 84.995 146.125 86.135 ;
        RECT 146.345 85.045 149.855 86.135 ;
        RECT 144.590 84.795 145.330 84.825 ;
        RECT 143.305 84.195 143.835 84.365 ;
        RECT 141.615 83.775 141.965 83.945 ;
        RECT 142.185 83.755 143.135 84.035 ;
        RECT 143.305 83.585 143.495 84.025 ;
        RECT 143.665 83.965 143.835 84.195 ;
        RECT 144.005 84.135 144.245 84.535 ;
        RECT 144.415 84.495 145.330 84.795 ;
        RECT 144.415 84.320 144.740 84.495 ;
        RECT 144.415 83.965 144.735 84.320 ;
        RECT 145.500 84.295 145.705 84.945 ;
        RECT 146.345 84.355 147.995 84.875 ;
        RECT 148.165 84.525 149.855 85.045 ;
        RECT 150.945 85.045 152.155 86.135 ;
        RECT 150.945 84.505 151.465 85.045 ;
        RECT 143.665 83.795 144.735 83.965 ;
        RECT 144.980 83.585 145.285 84.045 ;
        RECT 145.455 83.765 145.705 84.295 ;
        RECT 145.875 83.585 146.125 84.340 ;
        RECT 146.345 83.585 149.855 84.355 ;
        RECT 151.635 84.335 152.155 84.875 ;
        RECT 150.945 83.585 152.155 84.335 ;
        RECT 91.060 83.415 152.240 83.585 ;
        RECT 91.145 82.665 92.355 83.415 ;
        RECT 92.525 82.870 97.870 83.415 ;
        RECT 98.045 82.870 103.390 83.415 ;
        RECT 103.565 82.870 108.910 83.415 ;
        RECT 91.145 82.125 91.665 82.665 ;
        RECT 91.835 81.955 92.355 82.495 ;
        RECT 94.110 82.040 94.450 82.870 ;
        RECT 91.145 80.865 92.355 81.955 ;
        RECT 95.930 81.300 96.280 82.550 ;
        RECT 99.630 82.040 99.970 82.870 ;
        RECT 101.450 81.300 101.800 82.550 ;
        RECT 105.150 82.040 105.490 82.870 ;
        RECT 109.085 82.645 112.595 83.415 ;
        RECT 106.970 81.300 107.320 82.550 ;
        RECT 109.085 82.125 110.735 82.645 ;
        RECT 113.725 82.595 113.955 83.415 ;
        RECT 114.125 82.615 114.455 83.245 ;
        RECT 110.905 81.955 112.595 82.475 ;
        RECT 113.705 82.175 114.035 82.425 ;
        RECT 114.205 82.015 114.455 82.615 ;
        RECT 114.625 82.595 114.835 83.415 ;
        RECT 115.065 82.740 115.325 83.245 ;
        RECT 115.505 83.035 115.835 83.415 ;
        RECT 116.015 82.865 116.185 83.245 ;
        RECT 92.525 80.865 97.870 81.300 ;
        RECT 98.045 80.865 103.390 81.300 ;
        RECT 103.565 80.865 108.910 81.300 ;
        RECT 109.085 80.865 112.595 81.955 ;
        RECT 113.725 80.865 113.955 82.005 ;
        RECT 114.125 81.035 114.455 82.015 ;
        RECT 114.625 80.865 114.835 82.005 ;
        RECT 115.065 81.940 115.235 82.740 ;
        RECT 115.520 82.695 116.185 82.865 ;
        RECT 115.520 82.440 115.690 82.695 ;
        RECT 116.905 82.690 117.195 83.415 ;
        RECT 117.365 82.765 117.625 83.245 ;
        RECT 117.795 82.875 118.045 83.415 ;
        RECT 115.405 82.110 115.690 82.440 ;
        RECT 115.925 82.145 116.255 82.515 ;
        RECT 115.520 81.965 115.690 82.110 ;
        RECT 115.065 81.035 115.335 81.940 ;
        RECT 115.520 81.795 116.185 81.965 ;
        RECT 115.505 80.865 115.835 81.625 ;
        RECT 116.015 81.035 116.185 81.795 ;
        RECT 116.905 80.865 117.195 82.030 ;
        RECT 117.365 81.735 117.535 82.765 ;
        RECT 118.215 82.710 118.435 83.195 ;
        RECT 117.705 82.115 117.935 82.510 ;
        RECT 118.105 82.285 118.435 82.710 ;
        RECT 118.605 83.035 119.495 83.205 ;
        RECT 118.605 82.310 118.775 83.035 ;
        RECT 120.750 82.905 120.990 83.415 ;
        RECT 121.170 82.905 121.450 83.235 ;
        RECT 121.680 82.905 121.895 83.415 ;
        RECT 118.945 82.480 119.495 82.865 ;
        RECT 118.605 82.240 119.495 82.310 ;
        RECT 118.600 82.215 119.495 82.240 ;
        RECT 118.590 82.200 119.495 82.215 ;
        RECT 118.585 82.185 119.495 82.200 ;
        RECT 118.575 82.180 119.495 82.185 ;
        RECT 118.570 82.170 119.495 82.180 ;
        RECT 120.645 82.175 121.000 82.735 ;
        RECT 118.565 82.160 119.495 82.170 ;
        RECT 118.555 82.155 119.495 82.160 ;
        RECT 118.545 82.145 119.495 82.155 ;
        RECT 118.535 82.140 119.495 82.145 ;
        RECT 118.535 82.135 118.870 82.140 ;
        RECT 118.520 82.130 118.870 82.135 ;
        RECT 118.505 82.120 118.870 82.130 ;
        RECT 118.480 82.115 118.870 82.120 ;
        RECT 117.705 82.110 118.870 82.115 ;
        RECT 117.705 82.075 118.840 82.110 ;
        RECT 117.705 82.050 118.805 82.075 ;
        RECT 117.705 82.020 118.775 82.050 ;
        RECT 117.705 81.990 118.755 82.020 ;
        RECT 117.705 81.960 118.735 81.990 ;
        RECT 117.705 81.950 118.665 81.960 ;
        RECT 117.705 81.940 118.640 81.950 ;
        RECT 117.705 81.925 118.620 81.940 ;
        RECT 117.705 81.910 118.600 81.925 ;
        RECT 117.810 81.900 118.595 81.910 ;
        RECT 117.810 81.865 118.580 81.900 ;
        RECT 117.365 81.035 117.640 81.735 ;
        RECT 117.810 81.615 118.565 81.865 ;
        RECT 118.735 81.545 119.065 81.790 ;
        RECT 119.235 81.690 119.495 82.140 ;
        RECT 121.170 82.005 121.340 82.905 ;
        RECT 121.510 82.175 121.775 82.735 ;
        RECT 122.065 82.675 122.680 83.245 ;
        RECT 122.890 82.865 123.145 83.155 ;
        RECT 123.315 83.035 123.645 83.415 ;
        RECT 122.890 82.695 123.640 82.865 ;
        RECT 122.025 82.005 122.195 82.505 ;
        RECT 120.770 81.835 122.195 82.005 ;
        RECT 120.770 81.660 121.160 81.835 ;
        RECT 118.880 81.520 119.065 81.545 ;
        RECT 118.880 81.420 119.495 81.520 ;
        RECT 117.810 80.865 118.065 81.410 ;
        RECT 118.235 81.035 118.715 81.375 ;
        RECT 118.890 80.865 119.495 81.420 ;
        RECT 121.645 80.865 121.975 81.665 ;
        RECT 122.365 81.655 122.680 82.675 ;
        RECT 122.890 81.875 123.240 82.525 ;
        RECT 123.410 81.705 123.640 82.695 ;
        RECT 122.145 81.035 122.680 81.655 ;
        RECT 122.890 81.535 123.640 81.705 ;
        RECT 122.890 81.035 123.145 81.535 ;
        RECT 123.315 80.865 123.645 81.365 ;
        RECT 123.815 81.035 123.985 83.155 ;
        RECT 124.345 83.055 124.675 83.415 ;
        RECT 124.845 83.025 125.340 83.195 ;
        RECT 125.545 83.025 126.400 83.195 ;
        RECT 124.215 81.835 124.675 82.885 ;
        RECT 124.155 81.050 124.480 81.835 ;
        RECT 124.845 81.665 125.015 83.025 ;
        RECT 125.185 82.115 125.535 82.735 ;
        RECT 125.705 82.515 126.060 82.735 ;
        RECT 125.705 81.925 125.875 82.515 ;
        RECT 126.230 82.315 126.400 83.025 ;
        RECT 127.275 82.955 127.605 83.415 ;
        RECT 127.815 83.055 128.165 83.225 ;
        RECT 126.605 82.485 127.395 82.735 ;
        RECT 127.815 82.665 128.075 83.055 ;
        RECT 128.385 82.965 129.335 83.245 ;
        RECT 129.505 82.975 129.695 83.415 ;
        RECT 129.865 83.035 130.935 83.205 ;
        RECT 127.565 82.315 127.735 82.495 ;
        RECT 124.845 81.495 125.240 81.665 ;
        RECT 125.410 81.535 125.875 81.925 ;
        RECT 126.045 82.145 127.735 82.315 ;
        RECT 125.070 81.365 125.240 81.495 ;
        RECT 126.045 81.365 126.215 82.145 ;
        RECT 127.905 81.975 128.075 82.665 ;
        RECT 126.575 81.805 128.075 81.975 ;
        RECT 128.265 82.005 128.475 82.795 ;
        RECT 128.645 82.175 128.995 82.795 ;
        RECT 129.165 82.185 129.335 82.965 ;
        RECT 129.865 82.805 130.035 83.035 ;
        RECT 129.505 82.635 130.035 82.805 ;
        RECT 129.505 82.355 129.725 82.635 ;
        RECT 130.205 82.465 130.445 82.865 ;
        RECT 129.165 82.015 129.570 82.185 ;
        RECT 129.905 82.095 130.445 82.465 ;
        RECT 130.615 82.680 130.935 83.035 ;
        RECT 131.180 82.955 131.485 83.415 ;
        RECT 131.655 82.705 131.905 83.235 ;
        RECT 130.615 82.505 130.940 82.680 ;
        RECT 130.615 82.205 131.530 82.505 ;
        RECT 130.790 82.175 131.530 82.205 ;
        RECT 128.265 81.845 128.940 82.005 ;
        RECT 129.400 81.925 129.570 82.015 ;
        RECT 128.265 81.835 129.230 81.845 ;
        RECT 127.905 81.665 128.075 81.805 ;
        RECT 124.650 80.865 124.900 81.325 ;
        RECT 125.070 81.035 125.320 81.365 ;
        RECT 125.535 81.035 126.215 81.365 ;
        RECT 126.385 81.465 127.460 81.635 ;
        RECT 127.905 81.495 128.465 81.665 ;
        RECT 128.770 81.545 129.230 81.835 ;
        RECT 129.400 81.755 130.620 81.925 ;
        RECT 126.385 81.125 126.555 81.465 ;
        RECT 126.790 80.865 127.120 81.295 ;
        RECT 127.290 81.125 127.460 81.465 ;
        RECT 127.755 80.865 128.125 81.325 ;
        RECT 128.295 81.035 128.465 81.495 ;
        RECT 129.400 81.375 129.570 81.755 ;
        RECT 130.790 81.585 130.960 82.175 ;
        RECT 131.700 82.055 131.905 82.705 ;
        RECT 132.075 82.660 132.325 83.415 ;
        RECT 133.005 82.785 133.345 83.245 ;
        RECT 133.515 82.955 133.685 83.415 ;
        RECT 134.315 82.980 134.675 83.245 ;
        RECT 134.320 82.975 134.675 82.980 ;
        RECT 134.325 82.965 134.675 82.975 ;
        RECT 134.330 82.960 134.675 82.965 ;
        RECT 134.335 82.950 134.675 82.960 ;
        RECT 134.915 82.955 135.085 83.415 ;
        RECT 134.340 82.945 134.675 82.950 ;
        RECT 134.350 82.935 134.675 82.945 ;
        RECT 134.360 82.925 134.675 82.935 ;
        RECT 133.855 82.785 134.185 82.865 ;
        RECT 133.005 82.595 134.185 82.785 ;
        RECT 134.375 82.785 134.675 82.925 ;
        RECT 134.375 82.595 135.085 82.785 ;
        RECT 128.700 81.035 129.570 81.375 ;
        RECT 130.160 81.415 130.960 81.585 ;
        RECT 129.740 80.865 129.990 81.325 ;
        RECT 130.160 81.125 130.330 81.415 ;
        RECT 130.510 80.865 130.840 81.245 ;
        RECT 131.180 80.865 131.485 82.005 ;
        RECT 131.655 81.175 131.905 82.055 ;
        RECT 133.005 82.225 133.335 82.425 ;
        RECT 133.645 82.405 133.975 82.425 ;
        RECT 133.525 82.225 133.975 82.405 ;
        RECT 132.075 80.865 132.325 82.005 ;
        RECT 133.005 81.885 133.235 82.225 ;
        RECT 133.015 80.865 133.345 81.585 ;
        RECT 133.525 81.110 133.740 82.225 ;
        RECT 134.145 82.195 134.615 82.425 ;
        RECT 134.800 82.025 135.085 82.595 ;
        RECT 135.255 82.470 135.595 83.245 ;
        RECT 133.935 81.810 135.085 82.025 ;
        RECT 133.935 81.035 134.265 81.810 ;
        RECT 134.435 80.865 135.145 81.640 ;
        RECT 135.315 81.035 135.595 82.470 ;
        RECT 135.765 82.645 137.435 83.415 ;
        RECT 135.765 82.125 136.515 82.645 ;
        RECT 138.125 82.595 138.335 83.415 ;
        RECT 138.505 82.615 138.835 83.245 ;
        RECT 136.685 81.955 137.435 82.475 ;
        RECT 138.505 82.015 138.755 82.615 ;
        RECT 139.005 82.595 139.235 83.415 ;
        RECT 139.445 82.645 142.035 83.415 ;
        RECT 142.665 82.690 142.955 83.415 ;
        RECT 138.925 82.175 139.255 82.425 ;
        RECT 139.445 82.125 140.655 82.645 ;
        RECT 143.185 82.595 143.395 83.415 ;
        RECT 143.565 82.615 143.895 83.245 ;
        RECT 135.765 80.865 137.435 81.955 ;
        RECT 138.125 80.865 138.335 82.005 ;
        RECT 138.505 81.035 138.835 82.015 ;
        RECT 139.005 80.865 139.235 82.005 ;
        RECT 140.825 81.955 142.035 82.475 ;
        RECT 139.445 80.865 142.035 81.955 ;
        RECT 142.665 80.865 142.955 82.030 ;
        RECT 143.565 82.015 143.815 82.615 ;
        RECT 144.065 82.595 144.295 83.415 ;
        RECT 144.505 82.870 149.850 83.415 ;
        RECT 143.985 82.175 144.315 82.425 ;
        RECT 146.090 82.040 146.430 82.870 ;
        RECT 150.945 82.665 152.155 83.415 ;
        RECT 143.185 80.865 143.395 82.005 ;
        RECT 143.565 81.035 143.895 82.015 ;
        RECT 144.065 80.865 144.295 82.005 ;
        RECT 147.910 81.300 148.260 82.550 ;
        RECT 150.945 81.955 151.465 82.495 ;
        RECT 151.635 82.125 152.155 82.665 ;
        RECT 144.505 80.865 149.850 81.300 ;
        RECT 150.945 80.865 152.155 81.955 ;
        RECT 91.060 80.695 152.240 80.865 ;
        RECT 91.145 79.605 92.355 80.695 ;
        RECT 92.525 80.260 97.870 80.695 ;
        RECT 98.045 80.260 103.390 80.695 ;
        RECT 91.145 78.895 91.665 79.435 ;
        RECT 91.835 79.065 92.355 79.605 ;
        RECT 91.145 78.145 92.355 78.895 ;
        RECT 94.110 78.690 94.450 79.520 ;
        RECT 95.930 79.010 96.280 80.260 ;
        RECT 99.630 78.690 99.970 79.520 ;
        RECT 101.450 79.010 101.800 80.260 ;
        RECT 104.025 79.530 104.315 80.695 ;
        RECT 104.485 80.260 109.830 80.695 ;
        RECT 92.525 78.145 97.870 78.690 ;
        RECT 98.045 78.145 103.390 78.690 ;
        RECT 104.025 78.145 104.315 78.870 ;
        RECT 106.070 78.690 106.410 79.520 ;
        RECT 107.890 79.010 108.240 80.260 ;
        RECT 110.930 80.025 111.185 80.525 ;
        RECT 111.355 80.195 111.685 80.695 ;
        RECT 110.930 79.855 111.680 80.025 ;
        RECT 110.930 79.035 111.280 79.685 ;
        RECT 111.450 78.865 111.680 79.855 ;
        RECT 110.930 78.695 111.680 78.865 ;
        RECT 104.485 78.145 109.830 78.690 ;
        RECT 110.930 78.405 111.185 78.695 ;
        RECT 111.355 78.145 111.685 78.525 ;
        RECT 111.855 78.405 112.025 80.525 ;
        RECT 112.195 79.725 112.520 80.510 ;
        RECT 112.690 80.235 112.940 80.695 ;
        RECT 113.110 80.195 113.360 80.525 ;
        RECT 113.575 80.195 114.255 80.525 ;
        RECT 113.110 80.065 113.280 80.195 ;
        RECT 112.885 79.895 113.280 80.065 ;
        RECT 112.255 78.675 112.715 79.725 ;
        RECT 112.885 78.535 113.055 79.895 ;
        RECT 113.450 79.635 113.915 80.025 ;
        RECT 113.225 78.825 113.575 79.445 ;
        RECT 113.745 79.045 113.915 79.635 ;
        RECT 114.085 79.415 114.255 80.195 ;
        RECT 114.425 80.095 114.595 80.435 ;
        RECT 114.830 80.265 115.160 80.695 ;
        RECT 115.330 80.095 115.500 80.435 ;
        RECT 115.795 80.235 116.165 80.695 ;
        RECT 114.425 79.925 115.500 80.095 ;
        RECT 116.335 80.065 116.505 80.525 ;
        RECT 116.740 80.185 117.610 80.525 ;
        RECT 117.780 80.235 118.030 80.695 ;
        RECT 115.945 79.895 116.505 80.065 ;
        RECT 115.945 79.755 116.115 79.895 ;
        RECT 114.615 79.585 116.115 79.755 ;
        RECT 116.810 79.725 117.270 80.015 ;
        RECT 114.085 79.245 115.775 79.415 ;
        RECT 113.745 78.825 114.100 79.045 ;
        RECT 114.270 78.535 114.440 79.245 ;
        RECT 114.645 78.825 115.435 79.075 ;
        RECT 115.605 79.065 115.775 79.245 ;
        RECT 115.945 78.895 116.115 79.585 ;
        RECT 112.385 78.145 112.715 78.505 ;
        RECT 112.885 78.365 113.380 78.535 ;
        RECT 113.585 78.365 114.440 78.535 ;
        RECT 115.315 78.145 115.645 78.605 ;
        RECT 115.855 78.505 116.115 78.895 ;
        RECT 116.305 79.715 117.270 79.725 ;
        RECT 117.440 79.805 117.610 80.185 ;
        RECT 118.200 80.145 118.370 80.435 ;
        RECT 118.550 80.315 118.880 80.695 ;
        RECT 118.200 79.975 119.000 80.145 ;
        RECT 116.305 79.555 116.980 79.715 ;
        RECT 117.440 79.635 118.660 79.805 ;
        RECT 116.305 78.765 116.515 79.555 ;
        RECT 117.440 79.545 117.610 79.635 ;
        RECT 116.685 78.765 117.035 79.385 ;
        RECT 117.205 79.375 117.610 79.545 ;
        RECT 117.205 78.595 117.375 79.375 ;
        RECT 117.545 78.925 117.765 79.205 ;
        RECT 117.945 79.095 118.485 79.465 ;
        RECT 118.830 79.385 119.000 79.975 ;
        RECT 119.220 79.555 119.525 80.695 ;
        RECT 119.695 79.505 119.945 80.385 ;
        RECT 120.115 79.555 120.365 80.695 ;
        RECT 121.505 80.140 122.110 80.695 ;
        RECT 122.285 80.185 122.765 80.525 ;
        RECT 122.935 80.150 123.190 80.695 ;
        RECT 121.505 80.040 122.120 80.140 ;
        RECT 121.935 80.015 122.120 80.040 ;
        RECT 118.830 79.355 119.570 79.385 ;
        RECT 117.545 78.755 118.075 78.925 ;
        RECT 115.855 78.335 116.205 78.505 ;
        RECT 116.425 78.315 117.375 78.595 ;
        RECT 117.545 78.145 117.735 78.585 ;
        RECT 117.905 78.525 118.075 78.755 ;
        RECT 118.245 78.695 118.485 79.095 ;
        RECT 118.655 79.055 119.570 79.355 ;
        RECT 118.655 78.880 118.980 79.055 ;
        RECT 118.655 78.525 118.975 78.880 ;
        RECT 119.740 78.855 119.945 79.505 ;
        RECT 121.505 79.420 121.765 79.870 ;
        RECT 121.935 79.770 122.265 80.015 ;
        RECT 122.435 79.695 123.190 79.945 ;
        RECT 123.360 79.825 123.635 80.525 ;
        RECT 124.725 80.185 125.025 80.695 ;
        RECT 125.195 80.015 125.525 80.525 ;
        RECT 125.695 80.185 126.325 80.695 ;
        RECT 126.905 80.185 127.285 80.355 ;
        RECT 127.455 80.185 127.755 80.695 ;
        RECT 127.115 80.015 127.285 80.185 ;
        RECT 122.420 79.660 123.190 79.695 ;
        RECT 122.405 79.650 123.190 79.660 ;
        RECT 122.400 79.635 123.295 79.650 ;
        RECT 122.380 79.620 123.295 79.635 ;
        RECT 122.360 79.610 123.295 79.620 ;
        RECT 122.335 79.600 123.295 79.610 ;
        RECT 122.265 79.570 123.295 79.600 ;
        RECT 122.245 79.540 123.295 79.570 ;
        RECT 122.225 79.510 123.295 79.540 ;
        RECT 122.195 79.485 123.295 79.510 ;
        RECT 122.160 79.450 123.295 79.485 ;
        RECT 122.130 79.445 123.295 79.450 ;
        RECT 122.130 79.440 122.520 79.445 ;
        RECT 122.130 79.430 122.495 79.440 ;
        RECT 122.130 79.425 122.480 79.430 ;
        RECT 122.130 79.420 122.465 79.425 ;
        RECT 121.505 79.415 122.465 79.420 ;
        RECT 121.505 79.405 122.455 79.415 ;
        RECT 121.505 79.400 122.445 79.405 ;
        RECT 121.505 79.390 122.435 79.400 ;
        RECT 121.505 79.380 122.430 79.390 ;
        RECT 121.505 79.375 122.425 79.380 ;
        RECT 121.505 79.360 122.415 79.375 ;
        RECT 121.505 79.345 122.410 79.360 ;
        RECT 121.505 79.320 122.400 79.345 ;
        RECT 121.505 79.250 122.395 79.320 ;
        RECT 117.905 78.355 118.975 78.525 ;
        RECT 119.220 78.145 119.525 78.605 ;
        RECT 119.695 78.325 119.945 78.855 ;
        RECT 120.115 78.145 120.365 78.900 ;
        RECT 121.505 78.695 122.055 79.080 ;
        RECT 122.225 78.525 122.395 79.250 ;
        RECT 121.505 78.355 122.395 78.525 ;
        RECT 122.565 78.850 122.895 79.275 ;
        RECT 123.065 79.050 123.295 79.445 ;
        RECT 122.565 78.365 122.785 78.850 ;
        RECT 123.465 78.795 123.635 79.825 ;
        RECT 122.955 78.145 123.205 78.685 ;
        RECT 123.375 78.315 123.635 78.795 ;
        RECT 124.725 79.845 126.945 80.015 ;
        RECT 124.725 78.885 124.895 79.845 ;
        RECT 125.065 79.505 126.605 79.675 ;
        RECT 125.065 79.055 125.310 79.505 ;
        RECT 125.570 79.135 126.265 79.335 ;
        RECT 126.435 79.305 126.605 79.505 ;
        RECT 126.775 79.645 126.945 79.845 ;
        RECT 127.115 79.815 127.775 80.015 ;
        RECT 126.775 79.475 127.435 79.645 ;
        RECT 126.435 79.135 127.035 79.305 ;
        RECT 127.265 79.055 127.435 79.475 ;
        RECT 124.725 78.340 125.190 78.885 ;
        RECT 125.695 78.145 125.865 78.965 ;
        RECT 126.035 78.885 126.945 78.965 ;
        RECT 127.605 78.885 127.775 79.815 ;
        RECT 127.985 79.555 128.215 80.695 ;
        RECT 128.385 79.545 128.715 80.525 ;
        RECT 128.885 79.555 129.095 80.695 ;
        RECT 127.965 79.135 128.295 79.385 ;
        RECT 126.035 78.795 127.285 78.885 ;
        RECT 126.035 78.315 126.365 78.795 ;
        RECT 126.775 78.715 127.285 78.795 ;
        RECT 126.535 78.145 126.885 78.535 ;
        RECT 127.055 78.315 127.285 78.715 ;
        RECT 127.455 78.405 127.775 78.885 ;
        RECT 127.985 78.145 128.215 78.965 ;
        RECT 128.465 78.945 128.715 79.545 ;
        RECT 129.785 79.530 130.075 80.695 ;
        RECT 131.170 80.305 131.505 80.525 ;
        RECT 132.510 80.315 132.865 80.695 ;
        RECT 131.170 79.685 131.425 80.305 ;
        RECT 131.675 80.145 131.905 80.185 ;
        RECT 133.035 80.145 133.285 80.525 ;
        RECT 131.675 79.945 133.285 80.145 ;
        RECT 131.675 79.855 131.860 79.945 ;
        RECT 132.450 79.935 133.285 79.945 ;
        RECT 133.535 79.915 133.785 80.695 ;
        RECT 133.955 79.845 134.215 80.525 ;
        RECT 132.015 79.745 132.345 79.775 ;
        RECT 132.015 79.685 133.815 79.745 ;
        RECT 131.170 79.575 133.875 79.685 ;
        RECT 131.170 79.515 132.345 79.575 ;
        RECT 133.675 79.540 133.875 79.575 ;
        RECT 131.165 79.135 131.655 79.335 ;
        RECT 131.845 79.135 132.320 79.345 ;
        RECT 128.385 78.315 128.715 78.945 ;
        RECT 128.885 78.145 129.095 78.965 ;
        RECT 129.785 78.145 130.075 78.870 ;
        RECT 131.170 78.145 131.625 78.910 ;
        RECT 132.100 78.735 132.320 79.135 ;
        RECT 132.565 79.135 132.895 79.345 ;
        RECT 132.565 78.735 132.775 79.135 ;
        RECT 133.065 79.100 133.475 79.405 ;
        RECT 133.705 78.965 133.875 79.540 ;
        RECT 133.605 78.845 133.875 78.965 ;
        RECT 133.030 78.800 133.875 78.845 ;
        RECT 133.030 78.675 133.785 78.800 ;
        RECT 133.030 78.525 133.200 78.675 ;
        RECT 134.045 78.645 134.215 79.845 ;
        RECT 131.900 78.315 133.200 78.525 ;
        RECT 133.455 78.145 133.785 78.505 ;
        RECT 133.955 78.315 134.215 78.645 ;
        RECT 134.390 79.745 134.655 80.515 ;
        RECT 134.825 79.975 135.155 80.695 ;
        RECT 135.345 80.155 135.605 80.515 ;
        RECT 135.775 80.325 136.105 80.695 ;
        RECT 136.275 80.155 136.535 80.515 ;
        RECT 135.345 79.925 136.535 80.155 ;
        RECT 137.105 79.745 137.395 80.515 ;
        RECT 137.605 80.260 142.950 80.695 ;
        RECT 134.390 78.325 134.725 79.745 ;
        RECT 134.900 79.565 137.395 79.745 ;
        RECT 134.900 78.875 135.125 79.565 ;
        RECT 135.325 79.055 135.605 79.385 ;
        RECT 135.785 79.055 136.360 79.385 ;
        RECT 136.540 79.055 136.975 79.385 ;
        RECT 137.155 79.055 137.425 79.385 ;
        RECT 134.900 78.685 137.385 78.875 ;
        RECT 139.190 78.690 139.530 79.520 ;
        RECT 141.010 79.010 141.360 80.260 ;
        RECT 143.125 79.555 143.395 80.525 ;
        RECT 143.605 79.895 143.885 80.695 ;
        RECT 144.065 80.145 145.260 80.475 ;
        RECT 144.390 79.725 144.810 79.975 ;
        RECT 143.565 79.555 144.810 79.725 ;
        RECT 143.125 78.820 143.295 79.555 ;
        RECT 143.565 79.385 143.735 79.555 ;
        RECT 145.035 79.385 145.205 79.945 ;
        RECT 145.455 79.555 145.710 80.695 ;
        RECT 145.885 79.605 149.395 80.695 ;
        RECT 149.565 79.605 150.775 80.695 ;
        RECT 143.505 79.055 143.735 79.385 ;
        RECT 144.465 79.055 145.205 79.385 ;
        RECT 145.375 79.135 145.710 79.385 ;
        RECT 143.565 78.885 143.735 79.055 ;
        RECT 144.955 78.965 145.205 79.055 ;
        RECT 134.905 78.145 135.650 78.515 ;
        RECT 136.215 78.325 136.470 78.685 ;
        RECT 136.650 78.145 136.980 78.515 ;
        RECT 137.160 78.325 137.385 78.685 ;
        RECT 137.605 78.145 142.950 78.690 ;
        RECT 143.125 78.475 143.395 78.820 ;
        RECT 143.565 78.715 144.305 78.885 ;
        RECT 144.955 78.795 145.690 78.965 ;
        RECT 143.585 78.145 143.965 78.545 ;
        RECT 144.135 78.365 144.305 78.715 ;
        RECT 144.475 78.145 145.210 78.625 ;
        RECT 145.380 78.325 145.690 78.795 ;
        RECT 145.885 78.915 147.535 79.435 ;
        RECT 147.705 79.085 149.395 79.605 ;
        RECT 145.885 78.145 149.395 78.915 ;
        RECT 149.565 78.895 150.085 79.435 ;
        RECT 150.255 79.065 150.775 79.605 ;
        RECT 150.945 79.605 152.155 80.695 ;
        RECT 150.945 79.065 151.465 79.605 ;
        RECT 151.635 78.895 152.155 79.435 ;
        RECT 149.565 78.145 150.775 78.895 ;
        RECT 150.945 78.145 152.155 78.895 ;
        RECT 91.060 77.975 152.240 78.145 ;
        RECT 91.145 77.225 92.355 77.975 ;
        RECT 92.525 77.430 97.870 77.975 ;
        RECT 98.045 77.430 103.390 77.975 ;
        RECT 91.145 76.685 91.665 77.225 ;
        RECT 91.835 76.515 92.355 77.055 ;
        RECT 94.110 76.600 94.450 77.430 ;
        RECT 91.145 75.425 92.355 76.515 ;
        RECT 95.930 75.860 96.280 77.110 ;
        RECT 99.630 76.600 99.970 77.430 ;
        RECT 103.565 77.205 107.075 77.975 ;
        RECT 107.245 77.225 108.455 77.975 ;
        RECT 108.625 77.300 108.885 77.805 ;
        RECT 109.065 77.595 109.395 77.975 ;
        RECT 109.575 77.425 109.745 77.805 ;
        RECT 110.005 77.430 115.350 77.975 ;
        RECT 101.450 75.860 101.800 77.110 ;
        RECT 103.565 76.685 105.215 77.205 ;
        RECT 105.385 76.515 107.075 77.035 ;
        RECT 107.245 76.685 107.765 77.225 ;
        RECT 107.935 76.515 108.455 77.055 ;
        RECT 92.525 75.425 97.870 75.860 ;
        RECT 98.045 75.425 103.390 75.860 ;
        RECT 103.565 75.425 107.075 76.515 ;
        RECT 107.245 75.425 108.455 76.515 ;
        RECT 108.625 76.500 108.795 77.300 ;
        RECT 109.080 77.255 109.745 77.425 ;
        RECT 109.080 77.000 109.250 77.255 ;
        RECT 108.965 76.670 109.250 77.000 ;
        RECT 109.485 76.705 109.815 77.075 ;
        RECT 109.080 76.525 109.250 76.670 ;
        RECT 111.590 76.600 111.930 77.430 ;
        RECT 115.525 77.225 116.735 77.975 ;
        RECT 116.905 77.250 117.195 77.975 ;
        RECT 117.365 77.225 118.575 77.975 ;
        RECT 118.745 77.595 119.635 77.765 ;
        RECT 108.625 75.595 108.895 76.500 ;
        RECT 109.080 76.355 109.745 76.525 ;
        RECT 109.065 75.425 109.395 76.185 ;
        RECT 109.575 75.595 109.745 76.355 ;
        RECT 113.410 75.860 113.760 77.110 ;
        RECT 115.525 76.685 116.045 77.225 ;
        RECT 116.215 76.515 116.735 77.055 ;
        RECT 117.365 76.685 117.885 77.225 ;
        RECT 110.005 75.425 115.350 75.860 ;
        RECT 115.525 75.425 116.735 76.515 ;
        RECT 116.905 75.425 117.195 76.590 ;
        RECT 118.055 76.515 118.575 77.055 ;
        RECT 118.745 77.040 119.295 77.425 ;
        RECT 119.465 76.870 119.635 77.595 ;
        RECT 117.365 75.425 118.575 76.515 ;
        RECT 118.745 76.800 119.635 76.870 ;
        RECT 119.805 77.270 120.025 77.755 ;
        RECT 120.195 77.435 120.445 77.975 ;
        RECT 120.615 77.325 120.875 77.805 ;
        RECT 119.805 76.845 120.135 77.270 ;
        RECT 118.745 76.775 119.640 76.800 ;
        RECT 118.745 76.760 119.650 76.775 ;
        RECT 118.745 76.745 119.655 76.760 ;
        RECT 118.745 76.740 119.665 76.745 ;
        RECT 118.745 76.730 119.670 76.740 ;
        RECT 118.745 76.720 119.675 76.730 ;
        RECT 118.745 76.715 119.685 76.720 ;
        RECT 118.745 76.705 119.695 76.715 ;
        RECT 118.745 76.700 119.705 76.705 ;
        RECT 118.745 76.250 119.005 76.700 ;
        RECT 119.370 76.695 119.705 76.700 ;
        RECT 119.370 76.690 119.720 76.695 ;
        RECT 119.370 76.680 119.735 76.690 ;
        RECT 119.370 76.675 119.760 76.680 ;
        RECT 120.305 76.675 120.535 77.070 ;
        RECT 119.370 76.670 120.535 76.675 ;
        RECT 119.400 76.635 120.535 76.670 ;
        RECT 119.435 76.610 120.535 76.635 ;
        RECT 119.465 76.580 120.535 76.610 ;
        RECT 119.485 76.550 120.535 76.580 ;
        RECT 119.505 76.520 120.535 76.550 ;
        RECT 119.575 76.510 120.535 76.520 ;
        RECT 119.600 76.500 120.535 76.510 ;
        RECT 119.620 76.485 120.535 76.500 ;
        RECT 119.640 76.470 120.535 76.485 ;
        RECT 119.645 76.460 120.430 76.470 ;
        RECT 119.660 76.425 120.430 76.460 ;
        RECT 119.175 76.105 119.505 76.350 ;
        RECT 119.675 76.175 120.430 76.425 ;
        RECT 120.705 76.295 120.875 77.325 ;
        RECT 121.105 77.155 121.315 77.975 ;
        RECT 121.485 77.175 121.815 77.805 ;
        RECT 121.485 76.575 121.735 77.175 ;
        RECT 121.985 77.155 122.215 77.975 ;
        RECT 122.425 77.430 127.770 77.975 ;
        RECT 121.905 76.735 122.235 76.985 ;
        RECT 124.010 76.600 124.350 77.430 ;
        RECT 127.945 77.205 131.455 77.975 ;
        RECT 131.625 77.255 131.965 77.765 ;
        RECT 119.175 76.080 119.360 76.105 ;
        RECT 118.745 75.980 119.360 76.080 ;
        RECT 118.745 75.425 119.350 75.980 ;
        RECT 119.525 75.595 120.005 75.935 ;
        RECT 120.175 75.425 120.430 75.970 ;
        RECT 120.600 75.595 120.875 76.295 ;
        RECT 121.105 75.425 121.315 76.565 ;
        RECT 121.485 75.595 121.815 76.575 ;
        RECT 121.985 75.425 122.215 76.565 ;
        RECT 125.830 75.860 126.180 77.110 ;
        RECT 127.945 76.685 129.595 77.205 ;
        RECT 129.765 76.515 131.455 77.035 ;
        RECT 122.425 75.425 127.770 75.860 ;
        RECT 127.945 75.425 131.455 76.515 ;
        RECT 131.625 75.855 131.885 77.255 ;
        RECT 132.135 77.175 132.405 77.975 ;
        RECT 132.060 76.735 132.390 76.985 ;
        RECT 132.585 76.735 132.865 77.705 ;
        RECT 133.045 76.735 133.345 77.705 ;
        RECT 133.525 76.735 133.875 77.700 ;
        RECT 134.095 77.475 134.590 77.805 ;
        RECT 132.075 76.565 132.390 76.735 ;
        RECT 134.095 76.565 134.265 77.475 ;
        RECT 132.075 76.395 134.265 76.565 ;
        RECT 131.625 75.595 131.965 75.855 ;
        RECT 132.135 75.425 132.465 76.225 ;
        RECT 132.930 75.595 133.180 76.395 ;
        RECT 133.365 75.425 133.695 76.145 ;
        RECT 133.915 75.595 134.165 76.395 ;
        RECT 134.435 75.985 134.675 77.295 ;
        RECT 134.335 75.425 134.670 75.805 ;
        RECT 134.845 75.595 135.125 77.695 ;
        RECT 135.355 77.515 135.525 77.975 ;
        RECT 135.795 77.585 137.045 77.765 ;
        RECT 136.180 77.345 136.545 77.415 ;
        RECT 135.295 77.165 136.545 77.345 ;
        RECT 136.715 77.365 137.045 77.585 ;
        RECT 137.215 77.535 137.385 77.975 ;
        RECT 137.555 77.365 137.895 77.780 ;
        RECT 136.715 77.195 137.895 77.365 ;
        RECT 138.065 77.205 140.655 77.975 ;
        RECT 140.830 77.445 141.120 77.795 ;
        RECT 141.315 77.615 141.645 77.975 ;
        RECT 141.815 77.445 142.045 77.750 ;
        RECT 140.830 77.275 142.045 77.445 ;
        RECT 135.295 76.565 135.570 77.165 ;
        RECT 135.740 76.735 136.095 76.985 ;
        RECT 136.290 76.955 136.755 76.985 ;
        RECT 136.285 76.785 136.755 76.955 ;
        RECT 136.290 76.735 136.755 76.785 ;
        RECT 136.925 76.735 137.255 76.985 ;
        RECT 137.430 76.785 137.895 76.985 ;
        RECT 137.075 76.615 137.255 76.735 ;
        RECT 138.065 76.685 139.275 77.205 ;
        RECT 142.235 77.105 142.405 77.670 ;
        RECT 142.665 77.250 142.955 77.975 ;
        RECT 135.295 76.355 136.905 76.565 ;
        RECT 137.075 76.445 137.405 76.615 ;
        RECT 136.495 76.255 136.905 76.355 ;
        RECT 135.315 75.425 136.100 76.185 ;
        RECT 136.495 75.595 136.880 76.255 ;
        RECT 137.205 75.655 137.405 76.445 ;
        RECT 137.575 75.425 137.895 76.605 ;
        RECT 139.445 76.515 140.655 77.035 ;
        RECT 140.890 76.955 141.150 77.065 ;
        RECT 140.885 76.785 141.150 76.955 ;
        RECT 140.890 76.735 141.150 76.785 ;
        RECT 141.330 76.735 141.715 77.065 ;
        RECT 141.885 76.935 142.405 77.105 ;
        RECT 143.125 77.235 143.590 77.780 ;
        RECT 138.065 75.425 140.655 76.515 ;
        RECT 140.830 75.425 141.150 76.565 ;
        RECT 141.330 75.685 141.525 76.735 ;
        RECT 141.885 76.555 142.055 76.935 ;
        RECT 141.705 76.275 142.055 76.555 ;
        RECT 142.245 76.405 142.490 76.765 ;
        RECT 141.705 75.595 142.035 76.275 ;
        RECT 142.235 75.425 142.490 76.225 ;
        RECT 142.665 75.425 142.955 76.590 ;
        RECT 143.125 76.275 143.295 77.235 ;
        RECT 144.095 77.155 144.265 77.975 ;
        RECT 144.435 77.325 144.765 77.805 ;
        RECT 144.935 77.585 145.285 77.975 ;
        RECT 145.455 77.405 145.685 77.805 ;
        RECT 145.175 77.325 145.685 77.405 ;
        RECT 144.435 77.235 145.685 77.325 ;
        RECT 145.855 77.235 146.175 77.715 ;
        RECT 144.435 77.155 145.345 77.235 ;
        RECT 143.465 76.615 143.710 77.065 ;
        RECT 143.970 76.785 144.665 76.985 ;
        RECT 144.835 76.815 145.435 76.985 ;
        RECT 144.835 76.615 145.005 76.815 ;
        RECT 145.665 76.645 145.835 77.065 ;
        RECT 143.465 76.445 145.005 76.615 ;
        RECT 145.175 76.475 145.835 76.645 ;
        RECT 145.175 76.275 145.345 76.475 ;
        RECT 146.005 76.305 146.175 77.235 ;
        RECT 146.385 77.155 146.615 77.975 ;
        RECT 146.785 77.175 147.115 77.805 ;
        RECT 146.365 76.735 146.695 76.985 ;
        RECT 146.865 76.575 147.115 77.175 ;
        RECT 147.285 77.155 147.495 77.975 ;
        RECT 147.725 77.205 150.315 77.975 ;
        RECT 150.945 77.225 152.155 77.975 ;
        RECT 147.725 76.685 148.935 77.205 ;
        RECT 143.125 76.105 145.345 76.275 ;
        RECT 145.515 76.105 146.175 76.305 ;
        RECT 143.125 75.425 143.425 75.935 ;
        RECT 143.595 75.595 143.925 76.105 ;
        RECT 145.515 75.935 145.685 76.105 ;
        RECT 144.095 75.425 144.725 75.935 ;
        RECT 145.305 75.765 145.685 75.935 ;
        RECT 145.855 75.425 146.155 75.935 ;
        RECT 146.385 75.425 146.615 76.565 ;
        RECT 146.785 75.595 147.115 76.575 ;
        RECT 147.285 75.425 147.495 76.565 ;
        RECT 149.105 76.515 150.315 77.035 ;
        RECT 147.725 75.425 150.315 76.515 ;
        RECT 150.945 76.515 151.465 77.055 ;
        RECT 151.635 76.685 152.155 77.225 ;
        RECT 150.945 75.425 152.155 76.515 ;
        RECT 91.060 75.255 152.240 75.425 ;
        RECT 91.145 74.165 92.355 75.255 ;
        RECT 92.525 74.820 97.870 75.255 ;
        RECT 98.045 74.820 103.390 75.255 ;
        RECT 91.145 73.455 91.665 73.995 ;
        RECT 91.835 73.625 92.355 74.165 ;
        RECT 91.145 72.705 92.355 73.455 ;
        RECT 94.110 73.250 94.450 74.080 ;
        RECT 95.930 73.570 96.280 74.820 ;
        RECT 99.630 73.250 99.970 74.080 ;
        RECT 101.450 73.570 101.800 74.820 ;
        RECT 104.025 74.090 104.315 75.255 ;
        RECT 104.490 74.585 104.745 75.085 ;
        RECT 104.915 74.755 105.245 75.255 ;
        RECT 104.490 74.415 105.240 74.585 ;
        RECT 104.490 73.595 104.840 74.245 ;
        RECT 92.525 72.705 97.870 73.250 ;
        RECT 98.045 72.705 103.390 73.250 ;
        RECT 104.025 72.705 104.315 73.430 ;
        RECT 105.010 73.425 105.240 74.415 ;
        RECT 104.490 73.255 105.240 73.425 ;
        RECT 104.490 72.965 104.745 73.255 ;
        RECT 104.915 72.705 105.245 73.085 ;
        RECT 105.415 72.965 105.585 75.085 ;
        RECT 105.755 74.285 106.080 75.070 ;
        RECT 106.250 74.795 106.500 75.255 ;
        RECT 106.670 74.755 106.920 75.085 ;
        RECT 107.135 74.755 107.815 75.085 ;
        RECT 106.670 74.625 106.840 74.755 ;
        RECT 106.445 74.455 106.840 74.625 ;
        RECT 105.815 73.235 106.275 74.285 ;
        RECT 106.445 73.095 106.615 74.455 ;
        RECT 107.010 74.195 107.475 74.585 ;
        RECT 106.785 73.385 107.135 74.005 ;
        RECT 107.305 73.605 107.475 74.195 ;
        RECT 107.645 73.975 107.815 74.755 ;
        RECT 107.985 74.655 108.155 74.995 ;
        RECT 108.390 74.825 108.720 75.255 ;
        RECT 108.890 74.655 109.060 74.995 ;
        RECT 109.355 74.795 109.725 75.255 ;
        RECT 107.985 74.485 109.060 74.655 ;
        RECT 109.895 74.625 110.065 75.085 ;
        RECT 110.300 74.745 111.170 75.085 ;
        RECT 111.340 74.795 111.590 75.255 ;
        RECT 109.505 74.455 110.065 74.625 ;
        RECT 109.505 74.315 109.675 74.455 ;
        RECT 108.175 74.145 109.675 74.315 ;
        RECT 110.370 74.285 110.830 74.575 ;
        RECT 107.645 73.805 109.335 73.975 ;
        RECT 107.305 73.385 107.660 73.605 ;
        RECT 107.830 73.095 108.000 73.805 ;
        RECT 108.205 73.385 108.995 73.635 ;
        RECT 109.165 73.625 109.335 73.805 ;
        RECT 109.505 73.455 109.675 74.145 ;
        RECT 105.945 72.705 106.275 73.065 ;
        RECT 106.445 72.925 106.940 73.095 ;
        RECT 107.145 72.925 108.000 73.095 ;
        RECT 108.875 72.705 109.205 73.165 ;
        RECT 109.415 73.065 109.675 73.455 ;
        RECT 109.865 74.275 110.830 74.285 ;
        RECT 111.000 74.365 111.170 74.745 ;
        RECT 111.760 74.705 111.930 74.995 ;
        RECT 112.110 74.875 112.440 75.255 ;
        RECT 111.760 74.535 112.560 74.705 ;
        RECT 109.865 74.115 110.540 74.275 ;
        RECT 111.000 74.195 112.220 74.365 ;
        RECT 109.865 73.325 110.075 74.115 ;
        RECT 111.000 74.105 111.170 74.195 ;
        RECT 110.245 73.325 110.595 73.945 ;
        RECT 110.765 73.935 111.170 74.105 ;
        RECT 110.765 73.155 110.935 73.935 ;
        RECT 111.105 73.485 111.325 73.765 ;
        RECT 111.505 73.655 112.045 74.025 ;
        RECT 112.390 73.915 112.560 74.535 ;
        RECT 112.735 74.195 112.905 75.255 ;
        RECT 113.115 74.245 113.405 75.085 ;
        RECT 113.575 74.415 113.745 75.255 ;
        RECT 113.955 74.245 114.205 75.085 ;
        RECT 114.415 74.415 114.585 75.255 ;
        RECT 115.065 74.745 115.365 75.255 ;
        RECT 115.535 74.575 115.865 75.085 ;
        RECT 116.035 74.745 116.665 75.255 ;
        RECT 117.245 74.745 117.625 74.915 ;
        RECT 117.795 74.745 118.095 75.255 ;
        RECT 117.455 74.575 117.625 74.745 ;
        RECT 115.065 74.405 117.285 74.575 ;
        RECT 113.115 74.075 114.840 74.245 ;
        RECT 111.105 73.315 111.635 73.485 ;
        RECT 109.415 72.895 109.765 73.065 ;
        RECT 109.985 72.875 110.935 73.155 ;
        RECT 111.105 72.705 111.295 73.145 ;
        RECT 111.465 73.085 111.635 73.315 ;
        RECT 111.805 73.255 112.045 73.655 ;
        RECT 112.215 73.905 112.560 73.915 ;
        RECT 112.215 73.695 114.245 73.905 ;
        RECT 112.215 73.440 112.540 73.695 ;
        RECT 114.430 73.525 114.840 74.075 ;
        RECT 112.215 73.085 112.535 73.440 ;
        RECT 111.465 72.915 112.535 73.085 ;
        RECT 112.735 72.705 112.905 73.515 ;
        RECT 113.075 73.355 114.840 73.525 ;
        RECT 115.065 73.445 115.235 74.405 ;
        RECT 115.405 74.065 116.945 74.235 ;
        RECT 115.405 73.615 115.650 74.065 ;
        RECT 115.910 73.695 116.605 73.895 ;
        RECT 116.775 73.865 116.945 74.065 ;
        RECT 117.115 74.205 117.285 74.405 ;
        RECT 117.455 74.375 118.115 74.575 ;
        RECT 117.115 74.035 117.775 74.205 ;
        RECT 116.775 73.695 117.375 73.865 ;
        RECT 117.605 73.615 117.775 74.035 ;
        RECT 113.075 72.875 113.405 73.355 ;
        RECT 113.575 72.705 113.745 73.175 ;
        RECT 113.915 72.875 114.245 73.355 ;
        RECT 114.415 72.705 114.585 73.175 ;
        RECT 115.065 72.900 115.530 73.445 ;
        RECT 116.035 72.705 116.205 73.525 ;
        RECT 116.375 73.445 117.285 73.525 ;
        RECT 117.945 73.445 118.115 74.375 ;
        RECT 118.285 74.165 119.495 75.255 ;
        RECT 116.375 73.355 117.625 73.445 ;
        RECT 116.375 72.875 116.705 73.355 ;
        RECT 117.115 73.275 117.625 73.355 ;
        RECT 116.875 72.705 117.225 73.095 ;
        RECT 117.395 72.875 117.625 73.275 ;
        RECT 117.795 72.965 118.115 73.445 ;
        RECT 118.285 73.455 118.805 73.995 ;
        RECT 118.975 73.625 119.495 74.165 ;
        RECT 119.675 74.195 120.005 75.045 ;
        RECT 118.285 72.705 119.495 73.455 ;
        RECT 119.675 73.430 119.865 74.195 ;
        RECT 120.175 74.115 120.425 75.255 ;
        RECT 120.615 74.615 120.865 75.035 ;
        RECT 121.095 74.785 121.425 75.255 ;
        RECT 121.655 74.615 121.905 75.035 ;
        RECT 120.615 74.445 121.905 74.615 ;
        RECT 122.085 74.615 122.415 75.045 ;
        RECT 122.085 74.445 122.540 74.615 ;
        RECT 120.605 73.945 120.820 74.275 ;
        RECT 120.035 73.615 120.345 73.945 ;
        RECT 120.515 73.615 120.820 73.945 ;
        RECT 120.995 73.615 121.280 74.275 ;
        RECT 121.475 73.615 121.740 74.275 ;
        RECT 121.955 73.615 122.200 74.275 ;
        RECT 120.175 73.445 120.345 73.615 ;
        RECT 122.370 73.445 122.540 74.445 ;
        RECT 122.885 74.165 125.475 75.255 ;
        RECT 119.675 72.920 120.005 73.430 ;
        RECT 120.175 73.275 122.540 73.445 ;
        RECT 122.885 73.475 124.095 73.995 ;
        RECT 124.265 73.645 125.475 74.165 ;
        RECT 126.140 74.465 126.675 75.085 ;
        RECT 120.175 72.705 120.505 73.105 ;
        RECT 121.555 72.935 121.885 73.275 ;
        RECT 122.055 72.705 122.385 73.105 ;
        RECT 122.885 72.705 125.475 73.475 ;
        RECT 126.140 73.445 126.455 74.465 ;
        RECT 126.845 74.455 127.175 75.255 ;
        RECT 127.660 74.285 128.050 74.460 ;
        RECT 126.625 74.115 128.050 74.285 ;
        RECT 128.405 74.165 129.615 75.255 ;
        RECT 126.625 73.615 126.795 74.115 ;
        RECT 126.140 72.875 126.755 73.445 ;
        RECT 127.045 73.385 127.310 73.945 ;
        RECT 127.480 73.215 127.650 74.115 ;
        RECT 127.820 73.385 128.175 73.945 ;
        RECT 128.405 73.455 128.925 73.995 ;
        RECT 129.095 73.625 129.615 74.165 ;
        RECT 129.785 74.090 130.075 75.255 ;
        RECT 130.710 74.305 130.975 75.075 ;
        RECT 131.145 74.535 131.475 75.255 ;
        RECT 131.665 74.715 131.925 75.075 ;
        RECT 132.095 74.885 132.425 75.255 ;
        RECT 132.595 74.715 132.855 75.075 ;
        RECT 131.665 74.485 132.855 74.715 ;
        RECT 133.425 74.305 133.715 75.075 ;
        RECT 133.925 74.820 139.270 75.255 ;
        RECT 126.925 72.705 127.140 73.215 ;
        RECT 127.370 72.885 127.650 73.215 ;
        RECT 127.830 72.705 128.070 73.215 ;
        RECT 128.405 72.705 129.615 73.455 ;
        RECT 129.785 72.705 130.075 73.430 ;
        RECT 130.710 72.885 131.045 74.305 ;
        RECT 131.220 74.125 133.715 74.305 ;
        RECT 131.220 73.435 131.445 74.125 ;
        RECT 131.645 73.615 131.925 73.945 ;
        RECT 132.105 73.615 132.680 73.945 ;
        RECT 132.860 73.615 133.295 73.945 ;
        RECT 133.475 73.615 133.745 73.945 ;
        RECT 131.220 73.245 133.705 73.435 ;
        RECT 135.510 73.250 135.850 74.080 ;
        RECT 137.330 73.570 137.680 74.820 ;
        RECT 139.445 74.165 140.655 75.255 ;
        RECT 139.445 73.455 139.965 73.995 ;
        RECT 140.135 73.625 140.655 74.165 ;
        RECT 140.885 74.115 141.095 75.255 ;
        RECT 141.265 74.105 141.595 75.085 ;
        RECT 141.765 74.115 141.995 75.255 ;
        RECT 142.665 74.115 142.945 75.255 ;
        RECT 143.115 74.105 143.445 75.085 ;
        RECT 143.615 74.115 143.875 75.255 ;
        RECT 144.045 74.115 144.385 75.085 ;
        RECT 144.555 74.115 144.725 75.255 ;
        RECT 144.995 74.455 145.245 75.255 ;
        RECT 145.890 74.285 146.220 75.085 ;
        RECT 146.520 74.455 146.850 75.255 ;
        RECT 147.020 74.285 147.350 75.085 ;
        RECT 144.915 74.115 147.350 74.285 ;
        RECT 147.725 74.165 150.315 75.255 ;
        RECT 131.225 72.705 131.970 73.075 ;
        RECT 132.535 72.885 132.790 73.245 ;
        RECT 132.970 72.705 133.300 73.075 ;
        RECT 133.480 72.885 133.705 73.245 ;
        RECT 133.925 72.705 139.270 73.250 ;
        RECT 139.445 72.705 140.655 73.455 ;
        RECT 140.885 72.705 141.095 73.525 ;
        RECT 141.265 73.505 141.515 74.105 ;
        RECT 141.685 73.695 142.015 73.945 ;
        RECT 142.675 73.675 143.010 73.945 ;
        RECT 141.265 72.875 141.595 73.505 ;
        RECT 141.765 72.705 141.995 73.525 ;
        RECT 143.180 73.505 143.350 74.105 ;
        RECT 143.520 73.695 143.855 73.945 ;
        RECT 144.045 73.555 144.220 74.115 ;
        RECT 144.915 73.865 145.085 74.115 ;
        RECT 144.390 73.695 145.085 73.865 ;
        RECT 145.260 73.695 145.680 73.895 ;
        RECT 145.850 73.695 146.180 73.895 ;
        RECT 146.350 73.695 146.680 73.895 ;
        RECT 144.045 73.505 144.275 73.555 ;
        RECT 142.665 72.705 142.975 73.505 ;
        RECT 143.180 72.875 143.875 73.505 ;
        RECT 144.045 72.875 144.385 73.505 ;
        RECT 144.555 72.705 144.805 73.505 ;
        RECT 144.995 73.355 146.220 73.525 ;
        RECT 144.995 72.875 145.325 73.355 ;
        RECT 145.495 72.705 145.720 73.165 ;
        RECT 145.890 72.875 146.220 73.355 ;
        RECT 146.850 73.485 147.020 74.115 ;
        RECT 147.205 73.695 147.555 73.945 ;
        RECT 146.850 72.875 147.350 73.485 ;
        RECT 147.725 73.475 148.935 73.995 ;
        RECT 149.105 73.645 150.315 74.165 ;
        RECT 150.945 74.165 152.155 75.255 ;
        RECT 150.945 73.625 151.465 74.165 ;
        RECT 147.725 72.705 150.315 73.475 ;
        RECT 151.635 73.455 152.155 73.995 ;
        RECT 150.945 72.705 152.155 73.455 ;
        RECT 91.060 72.535 152.240 72.705 ;
        RECT 23.400 71.850 23.830 72.300 ;
        RECT 32.795 71.800 33.470 72.475 ;
        RECT 91.145 71.785 92.355 72.535 ;
        RECT 92.525 71.990 97.870 72.535 ;
        RECT 98.045 71.990 103.390 72.535 ;
        RECT 91.145 71.245 91.665 71.785 ;
        RECT 23.480 71.105 23.830 71.215 ;
        RECT 22.330 70.935 23.830 71.105 ;
        RECT 21.890 69.810 22.060 70.370 ;
        RECT 19.055 69.640 22.060 69.810 ;
        RECT 19.055 69.630 20.865 69.640 ;
        RECT 19.055 67.875 19.425 69.630 ;
        RECT 21.890 69.330 22.060 69.640 ;
        RECT 21.890 68.120 22.060 68.700 ;
        RECT 21.135 67.940 22.060 68.120 ;
        RECT 18.850 66.960 19.580 67.875 ;
        RECT 21.135 67.385 21.330 67.940 ;
        RECT 21.890 67.660 22.060 67.940 ;
        RECT 19.990 67.225 20.500 67.310 ;
        RECT 21.025 67.225 21.545 67.385 ;
        RECT 19.990 67.015 21.545 67.225 ;
        RECT 22.330 67.335 22.500 70.935 ;
        RECT 23.480 70.855 23.830 70.935 ;
        RECT 24.750 70.855 26.790 71.025 ;
        RECT 23.575 67.335 23.935 67.460 ;
        RECT 22.330 67.155 23.935 67.335 ;
        RECT 23.575 67.100 23.935 67.155 ;
        RECT 19.070 64.485 19.420 66.960 ;
        RECT 19.990 66.940 20.500 67.015 ;
        RECT 21.025 66.875 21.545 67.015 ;
        RECT 22.995 66.880 23.325 66.935 ;
        RECT 21.140 66.135 21.325 66.875 ;
        RECT 22.340 66.700 23.325 66.880 ;
        RECT 24.310 66.760 24.480 70.650 ;
        RECT 24.750 67.660 24.920 70.855 ;
        RECT 21.900 66.135 22.070 66.410 ;
        RECT 21.140 65.950 22.070 66.135 ;
        RECT 21.900 65.370 22.070 65.950 ;
        RECT 21.900 64.485 22.070 64.740 ;
        RECT 19.070 64.260 22.070 64.485 ;
        RECT 19.070 63.720 19.415 64.260 ;
        RECT 18.930 63.285 19.550 63.720 ;
        RECT 21.900 63.700 22.070 64.260 ;
        RECT 22.340 63.740 22.510 66.700 ;
        RECT 22.995 66.515 23.325 66.700 ;
        RECT 23.980 66.590 24.480 66.760 ;
        RECT 25.190 66.760 25.360 70.650 ;
        RECT 26.180 67.285 26.350 69.960 ;
        RECT 26.620 69.400 26.790 70.855 ;
        RECT 28.395 71.015 30.250 71.185 ;
        RECT 91.835 71.075 92.355 71.615 ;
        RECT 94.110 71.160 94.450 71.990 ;
        RECT 27.400 69.580 28.085 70.140 ;
        RECT 26.620 69.230 27.180 69.400 ;
        RECT 26.620 68.920 26.790 69.230 ;
        RECT 26.620 67.710 26.790 68.290 ;
        RECT 27.310 67.710 27.900 67.900 ;
        RECT 26.620 67.530 27.900 67.710 ;
        RECT 26.175 66.850 26.355 67.285 ;
        RECT 26.620 67.250 26.790 67.530 ;
        RECT 27.310 67.270 27.900 67.530 ;
        RECT 25.190 66.590 25.680 66.760 ;
        RECT 26.175 66.670 27.175 66.850 ;
        RECT 22.340 63.100 22.515 63.740 ;
        RECT 22.765 63.100 23.100 63.190 ;
        RECT 22.340 62.925 23.100 63.100 ;
        RECT 22.765 62.845 23.100 62.925 ;
        RECT 21.415 62.060 21.845 62.240 ;
        RECT 23.540 62.060 23.710 66.370 ;
        RECT 23.980 63.380 24.150 66.590 ;
        RECT 24.420 63.380 24.590 66.370 ;
        RECT 24.210 62.580 24.580 62.985 ;
        RECT 21.415 61.890 23.710 62.060 ;
        RECT 21.415 61.730 21.845 61.890 ;
        RECT 24.300 61.585 24.475 62.580 ;
        RECT 24.200 61.150 24.610 61.585 ;
        RECT 25.070 59.755 25.240 66.370 ;
        RECT 25.510 63.380 25.680 66.590 ;
        RECT 24.890 59.335 25.425 59.755 ;
        RECT 6.030 58.825 6.380 58.830 ;
        RECT 6.030 57.510 8.240 58.825 ;
        RECT 25.950 58.165 26.120 66.370 ;
        RECT 26.560 65.135 26.730 66.370 ;
        RECT 27.000 66.090 27.170 66.670 ;
        RECT 27.000 65.910 27.500 66.090 ;
        RECT 27.000 65.330 27.170 65.910 ;
        RECT 28.395 65.135 28.565 71.015 ;
        RECT 29.640 66.760 29.810 70.650 ;
        RECT 30.080 67.660 30.250 71.015 ;
        RECT 31.235 70.925 31.565 71.010 ;
        RECT 31.235 70.755 32.360 70.925 ;
        RECT 31.235 70.680 31.565 70.755 ;
        RECT 29.310 66.590 29.810 66.760 ;
        RECT 30.520 66.760 30.690 70.650 ;
        RECT 31.035 69.400 31.405 69.495 ;
        RECT 31.750 69.400 31.920 69.960 ;
        RECT 31.035 69.230 31.920 69.400 ;
        RECT 31.035 69.155 31.405 69.230 ;
        RECT 31.750 68.920 31.920 69.230 ;
        RECT 31.750 67.710 31.920 68.290 ;
        RECT 31.420 67.530 31.920 67.710 ;
        RECT 31.750 66.935 31.920 67.530 ;
        RECT 32.190 67.250 32.360 70.755 ;
        RECT 34.260 70.140 34.630 70.450 ;
        RECT 30.520 66.590 31.010 66.760 ;
        RECT 31.665 66.660 32.005 66.935 ;
        RECT 26.560 64.965 28.565 65.135 ;
        RECT 26.560 63.660 26.730 64.965 ;
        RECT 27.000 64.390 27.170 64.700 ;
        RECT 27.000 64.220 27.560 64.390 ;
        RECT 27.000 63.660 27.170 64.220 ;
        RECT 27.550 63.225 28.240 63.780 ;
        RECT 28.870 59.605 29.040 66.370 ;
        RECT 29.310 63.380 29.480 66.590 ;
        RECT 29.750 63.395 29.920 66.370 ;
        RECT 28.685 59.095 29.310 59.605 ;
        RECT 29.750 59.570 29.925 63.395 ;
        RECT 30.400 61.770 30.570 66.370 ;
        RECT 30.840 63.380 31.010 66.590 ;
        RECT 31.280 62.650 31.450 66.370 ;
        RECT 31.750 66.030 31.920 66.660 ;
        RECT 32.800 66.630 32.970 69.960 ;
        RECT 33.240 69.400 33.410 69.960 ;
        RECT 34.310 69.835 34.585 70.140 ;
        RECT 91.145 69.985 92.355 71.075 ;
        RECT 95.930 70.420 96.280 71.670 ;
        RECT 99.630 71.160 99.970 71.990 ;
        RECT 103.565 71.765 107.075 72.535 ;
        RECT 107.245 71.785 108.455 72.535 ;
        RECT 101.450 70.420 101.800 71.670 ;
        RECT 103.565 71.245 105.215 71.765 ;
        RECT 105.385 71.075 107.075 71.595 ;
        RECT 107.245 71.245 107.765 71.785 ;
        RECT 108.665 71.715 108.895 72.535 ;
        RECT 109.065 71.735 109.395 72.365 ;
        RECT 107.935 71.075 108.455 71.615 ;
        RECT 108.645 71.295 108.975 71.545 ;
        RECT 109.145 71.135 109.395 71.735 ;
        RECT 109.565 71.715 109.775 72.535 ;
        RECT 110.005 71.765 113.515 72.535 ;
        RECT 113.685 71.785 114.895 72.535 ;
        RECT 115.090 72.145 115.420 72.535 ;
        RECT 115.590 71.975 115.815 72.355 ;
        RECT 110.005 71.245 111.655 71.765 ;
        RECT 92.525 69.985 97.870 70.420 ;
        RECT 98.045 69.985 103.390 70.420 ;
        RECT 103.565 69.985 107.075 71.075 ;
        RECT 107.245 69.985 108.455 71.075 ;
        RECT 108.665 69.985 108.895 71.125 ;
        RECT 109.065 70.155 109.395 71.135 ;
        RECT 109.565 69.985 109.775 71.125 ;
        RECT 111.825 71.075 113.515 71.595 ;
        RECT 113.685 71.245 114.205 71.785 ;
        RECT 114.375 71.075 114.895 71.615 ;
        RECT 115.075 71.295 115.315 71.945 ;
        RECT 115.485 71.795 115.815 71.975 ;
        RECT 115.485 71.125 115.660 71.795 ;
        RECT 116.015 71.625 116.245 72.245 ;
        RECT 116.425 71.805 116.725 72.535 ;
        RECT 116.905 71.810 117.195 72.535 ;
        RECT 117.385 71.845 117.625 72.365 ;
        RECT 117.795 72.040 118.190 72.535 ;
        RECT 118.755 72.205 118.925 72.350 ;
        RECT 118.550 72.010 118.925 72.205 ;
        RECT 115.830 71.295 116.245 71.625 ;
        RECT 116.425 71.295 116.720 71.625 ;
        RECT 110.005 69.985 113.515 71.075 ;
        RECT 113.685 69.985 114.895 71.075 ;
        RECT 115.075 70.935 115.660 71.125 ;
        RECT 115.075 70.165 115.350 70.935 ;
        RECT 115.830 70.765 116.725 71.095 ;
        RECT 115.520 70.595 116.725 70.765 ;
        RECT 115.520 70.165 115.850 70.595 ;
        RECT 116.020 69.985 116.215 70.425 ;
        RECT 116.395 70.165 116.725 70.595 ;
        RECT 116.905 69.985 117.195 71.150 ;
        RECT 117.385 71.040 117.560 71.845 ;
        RECT 118.550 71.675 118.720 72.010 ;
        RECT 119.205 71.965 119.445 72.340 ;
        RECT 119.615 72.030 119.950 72.535 ;
        RECT 119.205 71.815 119.425 71.965 ;
        RECT 117.735 71.315 118.720 71.675 ;
        RECT 118.890 71.485 119.425 71.815 ;
        RECT 117.735 71.295 119.020 71.315 ;
        RECT 118.160 71.145 119.020 71.295 ;
        RECT 117.385 70.255 117.690 71.040 ;
        RECT 117.865 70.665 118.560 70.975 ;
        RECT 117.870 69.985 118.555 70.455 ;
        RECT 118.735 70.200 119.020 71.145 ;
        RECT 119.190 70.835 119.425 71.485 ;
        RECT 119.595 71.005 119.895 71.855 ;
        RECT 120.125 71.785 121.335 72.535 ;
        RECT 121.620 71.905 121.905 72.365 ;
        RECT 122.075 72.075 122.345 72.535 ;
        RECT 120.125 71.245 120.645 71.785 ;
        RECT 121.620 71.735 122.575 71.905 ;
        RECT 120.815 71.075 121.335 71.615 ;
        RECT 119.190 70.605 119.865 70.835 ;
        RECT 119.195 69.985 119.525 70.435 ;
        RECT 119.695 70.175 119.865 70.605 ;
        RECT 120.125 69.985 121.335 71.075 ;
        RECT 121.505 71.005 122.195 71.565 ;
        RECT 122.365 70.835 122.575 71.735 ;
        RECT 121.620 70.615 122.575 70.835 ;
        RECT 122.745 71.565 123.145 72.365 ;
        RECT 123.335 71.905 123.615 72.365 ;
        RECT 124.135 72.075 124.460 72.535 ;
        RECT 123.335 71.735 124.460 71.905 ;
        RECT 124.630 71.795 125.015 72.365 ;
        RECT 124.010 71.625 124.460 71.735 ;
        RECT 122.745 71.005 123.840 71.565 ;
        RECT 124.010 71.295 124.565 71.625 ;
        RECT 121.620 70.155 121.905 70.615 ;
        RECT 122.075 69.985 122.345 70.445 ;
        RECT 122.745 70.155 123.145 71.005 ;
        RECT 124.010 70.835 124.460 71.295 ;
        RECT 124.735 71.125 125.015 71.795 ;
        RECT 125.195 71.725 125.465 72.535 ;
        RECT 125.635 71.725 125.965 72.365 ;
        RECT 126.135 71.725 126.375 72.535 ;
        RECT 126.590 72.145 126.920 72.535 ;
        RECT 127.090 71.975 127.315 72.355 ;
        RECT 125.185 71.295 125.535 71.545 ;
        RECT 125.705 71.125 125.875 71.725 ;
        RECT 126.045 71.295 126.395 71.545 ;
        RECT 126.575 71.295 126.815 71.945 ;
        RECT 126.985 71.795 127.315 71.975 ;
        RECT 126.985 71.125 127.160 71.795 ;
        RECT 127.515 71.625 127.745 72.245 ;
        RECT 127.925 71.805 128.225 72.535 ;
        RECT 128.405 71.765 131.915 72.535 ;
        RECT 132.085 71.785 133.295 72.535 ;
        RECT 133.465 71.795 133.905 72.355 ;
        RECT 134.075 71.795 134.525 72.535 ;
        RECT 134.695 71.965 134.865 72.365 ;
        RECT 135.035 72.135 135.455 72.535 ;
        RECT 135.625 71.965 135.855 72.365 ;
        RECT 134.695 71.795 135.855 71.965 ;
        RECT 136.025 71.795 136.515 72.365 ;
        RECT 127.330 71.295 127.745 71.625 ;
        RECT 127.925 71.295 128.220 71.625 ;
        RECT 128.405 71.245 130.055 71.765 ;
        RECT 123.335 70.615 124.460 70.835 ;
        RECT 123.335 70.155 123.615 70.615 ;
        RECT 124.135 69.985 124.460 70.445 ;
        RECT 124.630 70.155 125.015 71.125 ;
        RECT 125.195 69.985 125.525 71.125 ;
        RECT 125.705 70.955 126.385 71.125 ;
        RECT 126.055 70.170 126.385 70.955 ;
        RECT 126.575 70.935 127.160 71.125 ;
        RECT 126.575 70.165 126.850 70.935 ;
        RECT 127.330 70.765 128.225 71.095 ;
        RECT 130.225 71.075 131.915 71.595 ;
        RECT 132.085 71.245 132.605 71.785 ;
        RECT 132.775 71.075 133.295 71.615 ;
        RECT 127.020 70.595 128.225 70.765 ;
        RECT 127.020 70.165 127.350 70.595 ;
        RECT 127.520 69.985 127.715 70.425 ;
        RECT 127.895 70.165 128.225 70.595 ;
        RECT 128.405 69.985 131.915 71.075 ;
        RECT 132.085 69.985 133.295 71.075 ;
        RECT 133.465 70.785 133.775 71.795 ;
        RECT 133.945 71.175 134.115 71.625 ;
        RECT 134.285 71.345 134.675 71.625 ;
        RECT 134.860 71.295 135.105 71.625 ;
        RECT 133.945 71.005 134.735 71.175 ;
        RECT 133.465 70.155 133.905 70.785 ;
        RECT 134.080 69.985 134.395 70.835 ;
        RECT 134.565 70.325 134.735 71.005 ;
        RECT 134.905 70.495 135.105 71.295 ;
        RECT 135.305 70.495 135.555 71.625 ;
        RECT 135.770 71.295 136.175 71.625 ;
        RECT 136.345 71.125 136.515 71.795 ;
        RECT 136.745 71.715 136.955 72.535 ;
        RECT 137.125 71.735 137.455 72.365 ;
        RECT 137.125 71.135 137.375 71.735 ;
        RECT 137.625 71.715 137.855 72.535 ;
        RECT 138.585 71.715 138.795 72.535 ;
        RECT 138.965 71.735 139.295 72.365 ;
        RECT 137.545 71.295 137.875 71.545 ;
        RECT 138.965 71.135 139.215 71.735 ;
        RECT 139.465 71.715 139.695 72.535 ;
        RECT 139.910 72.030 140.245 72.535 ;
        RECT 140.415 71.965 140.655 72.340 ;
        RECT 140.935 72.205 141.105 72.350 ;
        RECT 140.935 72.010 141.310 72.205 ;
        RECT 141.670 72.040 142.065 72.535 ;
        RECT 139.385 71.295 139.715 71.545 ;
        RECT 135.745 70.955 136.515 71.125 ;
        RECT 135.745 70.325 135.995 70.955 ;
        RECT 134.565 70.155 135.995 70.325 ;
        RECT 136.175 69.985 136.505 70.785 ;
        RECT 136.745 69.985 136.955 71.125 ;
        RECT 137.125 70.155 137.455 71.135 ;
        RECT 137.625 69.985 137.855 71.125 ;
        RECT 138.585 69.985 138.795 71.125 ;
        RECT 138.965 70.155 139.295 71.135 ;
        RECT 139.465 69.985 139.695 71.125 ;
        RECT 139.965 71.005 140.265 71.855 ;
        RECT 140.435 71.815 140.655 71.965 ;
        RECT 140.435 71.485 140.970 71.815 ;
        RECT 141.140 71.675 141.310 72.010 ;
        RECT 142.235 71.845 142.475 72.365 ;
        RECT 140.435 70.835 140.670 71.485 ;
        RECT 141.140 71.315 142.125 71.675 ;
        RECT 139.995 70.605 140.670 70.835 ;
        RECT 140.840 71.295 142.125 71.315 ;
        RECT 140.840 71.145 141.700 71.295 ;
        RECT 139.995 70.175 140.165 70.605 ;
        RECT 140.335 69.985 140.665 70.435 ;
        RECT 140.840 70.200 141.125 71.145 ;
        RECT 142.300 71.040 142.475 71.845 ;
        RECT 142.665 71.810 142.955 72.535 ;
        RECT 143.125 71.715 143.385 72.535 ;
        RECT 143.555 71.715 143.885 72.135 ;
        RECT 144.065 72.050 144.855 72.315 ;
        RECT 143.635 71.625 143.885 71.715 ;
        RECT 141.300 70.665 141.995 70.975 ;
        RECT 141.305 69.985 141.990 70.455 ;
        RECT 142.170 70.255 142.475 71.040 ;
        RECT 142.665 69.985 142.955 71.150 ;
        RECT 143.125 70.665 143.465 71.545 ;
        RECT 143.635 71.375 144.430 71.625 ;
        RECT 143.125 69.985 143.385 70.495 ;
        RECT 143.635 70.155 143.805 71.375 ;
        RECT 144.600 71.195 144.855 72.050 ;
        RECT 145.025 71.895 145.225 72.315 ;
        RECT 145.415 72.075 145.745 72.535 ;
        RECT 145.025 71.375 145.435 71.895 ;
        RECT 145.915 71.885 146.175 72.365 ;
        RECT 145.605 71.195 145.835 71.625 ;
        RECT 144.045 71.025 145.835 71.195 ;
        RECT 144.045 70.660 144.295 71.025 ;
        RECT 144.465 70.665 144.795 70.855 ;
        RECT 145.015 70.730 145.730 71.025 ;
        RECT 146.005 70.855 146.175 71.885 ;
        RECT 144.465 70.490 144.660 70.665 ;
        RECT 144.045 69.985 144.660 70.490 ;
        RECT 144.830 70.155 145.305 70.495 ;
        RECT 145.475 69.985 145.690 70.530 ;
        RECT 145.900 70.155 146.175 70.855 ;
        RECT 146.345 71.795 146.605 72.365 ;
        RECT 146.775 72.135 147.160 72.535 ;
        RECT 147.330 71.965 147.585 72.365 ;
        RECT 146.775 71.795 147.585 71.965 ;
        RECT 147.775 71.795 148.020 72.365 ;
        RECT 148.190 72.135 148.575 72.535 ;
        RECT 148.745 71.965 149.000 72.365 ;
        RECT 148.190 71.795 149.000 71.965 ;
        RECT 149.190 71.795 149.615 72.365 ;
        RECT 149.785 72.135 150.170 72.535 ;
        RECT 150.340 71.965 150.775 72.365 ;
        RECT 149.785 71.795 150.775 71.965 ;
        RECT 146.345 71.125 146.530 71.795 ;
        RECT 146.775 71.625 147.125 71.795 ;
        RECT 147.775 71.625 147.945 71.795 ;
        RECT 148.190 71.625 148.540 71.795 ;
        RECT 149.190 71.625 149.540 71.795 ;
        RECT 149.785 71.625 150.120 71.795 ;
        RECT 150.945 71.785 152.155 72.535 ;
        RECT 146.700 71.295 147.125 71.625 ;
        RECT 146.345 70.155 146.605 71.125 ;
        RECT 146.775 70.775 147.125 71.295 ;
        RECT 147.295 71.125 147.945 71.625 ;
        RECT 148.115 71.295 148.540 71.625 ;
        RECT 147.295 70.945 148.020 71.125 ;
        RECT 146.775 70.580 147.585 70.775 ;
        RECT 146.775 69.985 147.160 70.410 ;
        RECT 147.330 70.155 147.585 70.580 ;
        RECT 147.775 70.155 148.020 70.945 ;
        RECT 148.190 70.775 148.540 71.295 ;
        RECT 148.710 71.125 149.540 71.625 ;
        RECT 149.710 71.295 150.120 71.625 ;
        RECT 148.710 70.945 149.615 71.125 ;
        RECT 148.190 70.580 149.020 70.775 ;
        RECT 148.190 69.985 148.575 70.410 ;
        RECT 148.745 70.155 149.020 70.580 ;
        RECT 149.190 70.155 149.615 70.945 ;
        RECT 149.785 70.750 150.120 71.295 ;
        RECT 150.290 70.920 150.775 71.625 ;
        RECT 150.945 71.075 151.465 71.615 ;
        RECT 151.635 71.245 152.155 71.785 ;
        RECT 149.785 70.580 150.775 70.750 ;
        RECT 149.785 69.985 150.170 70.410 ;
        RECT 150.340 70.155 150.775 70.580 ;
        RECT 150.945 69.985 152.155 71.075 ;
        RECT 34.080 69.455 34.810 69.835 ;
        RECT 91.060 69.815 152.240 69.985 ;
        RECT 34.080 69.400 35.445 69.455 ;
        RECT 33.240 69.285 35.445 69.400 ;
        RECT 33.240 69.230 34.810 69.285 ;
        RECT 33.240 68.920 33.410 69.230 ;
        RECT 34.080 68.885 34.810 69.230 ;
        RECT 33.240 67.710 33.410 68.290 ;
        RECT 33.755 67.710 34.255 67.865 ;
        RECT 33.240 67.530 34.255 67.710 ;
        RECT 33.240 67.250 33.410 67.530 ;
        RECT 33.755 67.350 34.255 67.530 ;
        RECT 33.940 66.985 34.110 67.350 ;
        RECT 33.840 66.655 34.250 66.985 ;
        RECT 32.095 66.030 32.265 66.310 ;
        RECT 31.750 65.850 32.265 66.030 ;
        RECT 32.095 65.270 32.265 65.850 ;
        RECT 31.630 65.000 31.960 65.080 ;
        RECT 32.535 65.000 32.705 66.310 ;
        RECT 31.630 64.830 32.705 65.000 ;
        RECT 31.630 64.750 31.960 64.830 ;
        RECT 32.095 64.330 32.265 64.640 ;
        RECT 31.705 64.160 32.265 64.330 ;
        RECT 31.040 62.385 31.455 62.650 ;
        RECT 31.705 62.305 31.875 64.160 ;
        RECT 32.095 63.600 32.265 64.160 ;
        RECT 32.535 63.600 32.705 64.830 ;
        RECT 33.145 62.780 33.315 66.310 ;
        RECT 33.585 66.030 33.755 66.310 ;
        RECT 33.940 66.030 34.110 66.655 ;
        RECT 33.585 65.850 34.110 66.030 ;
        RECT 35.275 65.975 35.445 69.285 ;
        RECT 91.145 68.725 92.355 69.815 ;
        RECT 92.525 69.380 97.870 69.815 ;
        RECT 91.145 68.015 91.665 68.555 ;
        RECT 91.835 68.185 92.355 68.725 ;
        RECT 91.145 67.265 92.355 68.015 ;
        RECT 94.110 67.810 94.450 68.640 ;
        RECT 95.930 68.130 96.280 69.380 ;
        RECT 98.045 68.725 100.635 69.815 ;
        RECT 98.045 68.035 99.255 68.555 ;
        RECT 99.425 68.205 100.635 68.725 ;
        RECT 101.265 68.740 101.535 69.645 ;
        RECT 101.705 69.055 102.035 69.815 ;
        RECT 102.215 68.885 102.385 69.645 ;
        RECT 92.525 67.265 97.870 67.810 ;
        RECT 98.045 67.265 100.635 68.035 ;
        RECT 101.265 67.940 101.435 68.740 ;
        RECT 101.720 68.715 102.385 68.885 ;
        RECT 102.645 68.725 103.855 69.815 ;
        RECT 101.720 68.570 101.890 68.715 ;
        RECT 101.605 68.240 101.890 68.570 ;
        RECT 101.720 67.985 101.890 68.240 ;
        RECT 102.125 68.165 102.455 68.535 ;
        RECT 102.645 68.015 103.165 68.555 ;
        RECT 103.335 68.185 103.855 68.725 ;
        RECT 104.025 68.650 104.315 69.815 ;
        RECT 104.485 69.380 109.830 69.815 ;
        RECT 101.265 67.435 101.525 67.940 ;
        RECT 101.720 67.815 102.385 67.985 ;
        RECT 101.705 67.265 102.035 67.645 ;
        RECT 102.215 67.435 102.385 67.815 ;
        RECT 102.645 67.265 103.855 68.015 ;
        RECT 104.025 67.265 104.315 67.990 ;
        RECT 106.070 67.810 106.410 68.640 ;
        RECT 107.890 68.130 108.240 69.380 ;
        RECT 110.930 69.145 111.185 69.645 ;
        RECT 111.355 69.315 111.685 69.815 ;
        RECT 110.930 68.975 111.680 69.145 ;
        RECT 110.930 68.155 111.280 68.805 ;
        RECT 111.450 67.985 111.680 68.975 ;
        RECT 110.930 67.815 111.680 67.985 ;
        RECT 104.485 67.265 109.830 67.810 ;
        RECT 110.930 67.525 111.185 67.815 ;
        RECT 111.355 67.265 111.685 67.645 ;
        RECT 111.855 67.525 112.025 69.645 ;
        RECT 112.195 68.845 112.520 69.630 ;
        RECT 112.690 69.355 112.940 69.815 ;
        RECT 113.110 69.315 113.360 69.645 ;
        RECT 113.575 69.315 114.255 69.645 ;
        RECT 113.110 69.185 113.280 69.315 ;
        RECT 112.885 69.015 113.280 69.185 ;
        RECT 112.255 67.795 112.715 68.845 ;
        RECT 112.885 67.655 113.055 69.015 ;
        RECT 113.450 68.755 113.915 69.145 ;
        RECT 113.225 67.945 113.575 68.565 ;
        RECT 113.745 68.165 113.915 68.755 ;
        RECT 114.085 68.535 114.255 69.315 ;
        RECT 114.425 69.215 114.595 69.555 ;
        RECT 114.830 69.385 115.160 69.815 ;
        RECT 115.330 69.215 115.500 69.555 ;
        RECT 115.795 69.355 116.165 69.815 ;
        RECT 114.425 69.045 115.500 69.215 ;
        RECT 116.335 69.185 116.505 69.645 ;
        RECT 116.740 69.305 117.610 69.645 ;
        RECT 117.780 69.355 118.030 69.815 ;
        RECT 115.945 69.015 116.505 69.185 ;
        RECT 115.945 68.875 116.115 69.015 ;
        RECT 114.615 68.705 116.115 68.875 ;
        RECT 116.810 68.845 117.270 69.135 ;
        RECT 114.085 68.365 115.775 68.535 ;
        RECT 113.745 67.945 114.100 68.165 ;
        RECT 114.270 67.655 114.440 68.365 ;
        RECT 114.645 67.945 115.435 68.195 ;
        RECT 115.605 68.185 115.775 68.365 ;
        RECT 115.945 68.015 116.115 68.705 ;
        RECT 112.385 67.265 112.715 67.625 ;
        RECT 112.885 67.485 113.380 67.655 ;
        RECT 113.585 67.485 114.440 67.655 ;
        RECT 115.315 67.265 115.645 67.725 ;
        RECT 115.855 67.625 116.115 68.015 ;
        RECT 116.305 68.835 117.270 68.845 ;
        RECT 117.440 68.925 117.610 69.305 ;
        RECT 118.200 69.265 118.370 69.555 ;
        RECT 118.550 69.435 118.880 69.815 ;
        RECT 118.200 69.095 119.000 69.265 ;
        RECT 116.305 68.675 116.980 68.835 ;
        RECT 117.440 68.755 118.660 68.925 ;
        RECT 116.305 67.885 116.515 68.675 ;
        RECT 117.440 68.665 117.610 68.755 ;
        RECT 116.685 67.885 117.035 68.505 ;
        RECT 117.205 68.495 117.610 68.665 ;
        RECT 117.205 67.715 117.375 68.495 ;
        RECT 117.545 68.045 117.765 68.325 ;
        RECT 117.945 68.215 118.485 68.585 ;
        RECT 118.830 68.505 119.000 69.095 ;
        RECT 119.220 68.675 119.525 69.815 ;
        RECT 119.695 68.625 119.945 69.505 ;
        RECT 120.115 68.675 120.365 69.815 ;
        RECT 120.585 69.095 121.045 69.645 ;
        RECT 121.235 69.095 121.565 69.815 ;
        RECT 118.830 68.475 119.570 68.505 ;
        RECT 117.545 67.875 118.075 68.045 ;
        RECT 115.855 67.455 116.205 67.625 ;
        RECT 116.425 67.435 117.375 67.715 ;
        RECT 117.545 67.265 117.735 67.705 ;
        RECT 117.905 67.645 118.075 67.875 ;
        RECT 118.245 67.815 118.485 68.215 ;
        RECT 118.655 68.175 119.570 68.475 ;
        RECT 118.655 68.000 118.980 68.175 ;
        RECT 118.655 67.645 118.975 68.000 ;
        RECT 119.740 67.975 119.945 68.625 ;
        RECT 117.905 67.475 118.975 67.645 ;
        RECT 119.220 67.265 119.525 67.725 ;
        RECT 119.695 67.445 119.945 67.975 ;
        RECT 120.115 67.265 120.365 68.020 ;
        RECT 120.585 67.725 120.835 69.095 ;
        RECT 121.765 68.925 122.065 69.475 ;
        RECT 122.235 69.145 122.515 69.815 ;
        RECT 122.885 69.380 128.230 69.815 ;
        RECT 121.125 68.755 122.065 68.925 ;
        RECT 121.125 68.505 121.295 68.755 ;
        RECT 122.435 68.505 122.700 68.865 ;
        RECT 121.005 68.175 121.295 68.505 ;
        RECT 121.465 68.255 121.805 68.505 ;
        RECT 122.025 68.255 122.700 68.505 ;
        RECT 121.125 68.085 121.295 68.175 ;
        RECT 121.125 67.895 122.515 68.085 ;
        RECT 120.585 67.435 121.145 67.725 ;
        RECT 121.315 67.265 121.565 67.725 ;
        RECT 122.185 67.535 122.515 67.895 ;
        RECT 124.470 67.810 124.810 68.640 ;
        RECT 126.290 68.130 126.640 69.380 ;
        RECT 128.405 68.725 129.615 69.815 ;
        RECT 128.405 68.015 128.925 68.555 ;
        RECT 129.095 68.185 129.615 68.725 ;
        RECT 129.785 68.650 130.075 69.815 ;
        RECT 130.245 68.725 131.915 69.815 ;
        RECT 132.175 69.195 132.345 69.625 ;
        RECT 132.515 69.365 132.845 69.815 ;
        RECT 132.175 68.965 132.850 69.195 ;
        RECT 130.245 68.035 130.995 68.555 ;
        RECT 131.165 68.205 131.915 68.725 ;
        RECT 122.885 67.265 128.230 67.810 ;
        RECT 128.405 67.265 129.615 68.015 ;
        RECT 129.785 67.265 130.075 67.990 ;
        RECT 130.245 67.265 131.915 68.035 ;
        RECT 132.145 67.945 132.445 68.795 ;
        RECT 132.615 68.315 132.850 68.965 ;
        RECT 133.020 68.655 133.305 69.600 ;
        RECT 133.485 69.345 134.170 69.815 ;
        RECT 133.480 68.825 134.175 69.135 ;
        RECT 134.350 68.760 134.655 69.545 ;
        RECT 133.020 68.505 133.880 68.655 ;
        RECT 133.020 68.485 134.305 68.505 ;
        RECT 132.615 67.985 133.150 68.315 ;
        RECT 133.320 68.125 134.305 68.485 ;
        RECT 132.615 67.835 132.835 67.985 ;
        RECT 132.090 67.265 132.425 67.770 ;
        RECT 132.595 67.460 132.835 67.835 ;
        RECT 133.320 67.790 133.490 68.125 ;
        RECT 134.480 67.955 134.655 68.760 ;
        RECT 134.850 68.675 135.105 69.815 ;
        RECT 135.300 69.265 136.495 69.595 ;
        RECT 135.355 68.505 135.525 69.065 ;
        RECT 135.750 68.845 136.170 69.095 ;
        RECT 136.675 69.015 136.955 69.815 ;
        RECT 135.750 68.675 136.995 68.845 ;
        RECT 137.165 68.675 137.435 69.645 ;
        RECT 137.610 68.675 137.865 69.815 ;
        RECT 138.060 69.265 139.255 69.595 ;
        RECT 136.825 68.505 136.995 68.675 ;
        RECT 134.850 68.255 135.185 68.505 ;
        RECT 135.355 68.175 136.095 68.505 ;
        RECT 136.825 68.175 137.055 68.505 ;
        RECT 135.355 68.085 135.605 68.175 ;
        RECT 133.115 67.595 133.490 67.790 ;
        RECT 133.115 67.450 133.285 67.595 ;
        RECT 133.850 67.265 134.245 67.760 ;
        RECT 134.415 67.435 134.655 67.955 ;
        RECT 134.870 67.915 135.605 68.085 ;
        RECT 136.825 68.005 136.995 68.175 ;
        RECT 134.870 67.445 135.180 67.915 ;
        RECT 136.255 67.835 136.995 68.005 ;
        RECT 137.265 67.940 137.435 68.675 ;
        RECT 138.115 68.505 138.285 69.065 ;
        RECT 138.510 68.845 138.930 69.095 ;
        RECT 139.435 69.015 139.715 69.815 ;
        RECT 138.510 68.675 139.755 68.845 ;
        RECT 139.925 68.675 140.195 69.645 ;
        RECT 140.365 68.725 142.035 69.815 ;
        RECT 139.585 68.505 139.755 68.675 ;
        RECT 137.610 68.255 137.945 68.505 ;
        RECT 138.115 68.175 138.855 68.505 ;
        RECT 139.585 68.175 139.815 68.505 ;
        RECT 138.115 68.085 138.365 68.175 ;
        RECT 135.350 67.265 136.085 67.745 ;
        RECT 136.255 67.485 136.425 67.835 ;
        RECT 136.595 67.265 136.975 67.665 ;
        RECT 137.165 67.595 137.435 67.940 ;
        RECT 137.630 67.915 138.365 68.085 ;
        RECT 139.585 68.005 139.755 68.175 ;
        RECT 137.630 67.445 137.940 67.915 ;
        RECT 139.015 67.835 139.755 68.005 ;
        RECT 140.025 67.940 140.195 68.675 ;
        RECT 138.110 67.265 138.845 67.745 ;
        RECT 139.015 67.485 139.185 67.835 ;
        RECT 139.355 67.265 139.735 67.665 ;
        RECT 139.925 67.595 140.195 67.940 ;
        RECT 140.365 68.035 141.115 68.555 ;
        RECT 141.285 68.205 142.035 68.725 ;
        RECT 142.755 68.805 142.925 69.645 ;
        RECT 143.095 69.475 144.265 69.645 ;
        RECT 143.095 68.975 143.425 69.475 ;
        RECT 143.935 69.435 144.265 69.475 ;
        RECT 144.455 69.395 144.810 69.815 ;
        RECT 143.595 69.215 143.825 69.305 ;
        RECT 144.980 69.215 145.230 69.645 ;
        RECT 143.595 68.975 145.230 69.215 ;
        RECT 145.400 69.055 145.730 69.815 ;
        RECT 145.900 68.975 146.155 69.645 ;
        RECT 142.755 68.635 145.815 68.805 ;
        RECT 142.670 68.255 143.020 68.465 ;
        RECT 143.190 68.255 143.635 68.455 ;
        RECT 143.805 68.255 144.280 68.455 ;
        RECT 140.365 67.265 142.035 68.035 ;
        RECT 142.755 67.915 143.820 68.085 ;
        RECT 142.755 67.435 142.925 67.915 ;
        RECT 143.095 67.265 143.425 67.745 ;
        RECT 143.650 67.685 143.820 67.915 ;
        RECT 144.000 67.855 144.280 68.255 ;
        RECT 144.550 68.255 144.880 68.455 ;
        RECT 145.050 68.255 145.415 68.455 ;
        RECT 144.550 67.855 144.835 68.255 ;
        RECT 145.645 68.085 145.815 68.635 ;
        RECT 145.015 67.915 145.815 68.085 ;
        RECT 145.015 67.685 145.185 67.915 ;
        RECT 145.985 67.845 146.155 68.975 ;
        RECT 145.970 67.765 146.155 67.845 ;
        RECT 143.650 67.435 145.185 67.685 ;
        RECT 145.355 67.265 145.685 67.745 ;
        RECT 145.900 67.435 146.155 67.765 ;
        RECT 146.345 68.675 146.615 69.645 ;
        RECT 146.825 69.015 147.105 69.815 ;
        RECT 147.285 69.265 148.480 69.595 ;
        RECT 147.610 68.845 148.030 69.095 ;
        RECT 146.785 68.675 148.030 68.845 ;
        RECT 146.345 68.625 146.575 68.675 ;
        RECT 146.345 67.940 146.515 68.625 ;
        RECT 146.785 68.505 146.955 68.675 ;
        RECT 148.255 68.505 148.425 69.065 ;
        RECT 148.675 68.675 148.930 69.815 ;
        RECT 149.105 68.725 150.775 69.815 ;
        RECT 146.725 68.175 146.955 68.505 ;
        RECT 147.685 68.175 148.425 68.505 ;
        RECT 148.595 68.255 148.930 68.505 ;
        RECT 146.785 68.005 146.955 68.175 ;
        RECT 148.175 68.085 148.425 68.175 ;
        RECT 146.345 67.595 146.615 67.940 ;
        RECT 146.785 67.835 147.525 68.005 ;
        RECT 148.175 67.915 148.910 68.085 ;
        RECT 146.805 67.265 147.185 67.665 ;
        RECT 147.355 67.485 147.525 67.835 ;
        RECT 147.695 67.265 148.430 67.745 ;
        RECT 148.600 67.445 148.910 67.915 ;
        RECT 149.105 68.035 149.855 68.555 ;
        RECT 150.025 68.205 150.775 68.725 ;
        RECT 150.945 68.725 152.155 69.815 ;
        RECT 150.945 68.185 151.465 68.725 ;
        RECT 149.105 67.265 150.775 68.035 ;
        RECT 151.635 68.015 152.155 68.555 ;
        RECT 150.945 67.265 152.155 68.015 ;
        RECT 91.060 67.095 152.240 67.265 ;
        RECT 91.145 66.345 92.355 67.095 ;
        RECT 92.525 66.550 97.870 67.095 ;
        RECT 33.585 65.270 33.755 65.850 ;
        RECT 35.135 65.595 35.590 65.975 ;
        RECT 91.145 65.805 91.665 66.345 ;
        RECT 91.835 65.635 92.355 66.175 ;
        RECT 94.110 65.720 94.450 66.550 ;
        RECT 98.510 66.545 98.765 66.835 ;
        RECT 98.935 66.715 99.265 67.095 ;
        RECT 98.510 66.375 99.260 66.545 ;
        RECT 33.585 64.330 33.755 64.640 ;
        RECT 34.430 64.585 34.980 65.080 ;
        RECT 34.455 64.580 34.835 64.585 ;
        RECT 35.275 64.330 35.445 65.595 ;
        RECT 91.145 64.545 92.355 65.635 ;
        RECT 95.930 64.980 96.280 66.230 ;
        RECT 98.510 65.555 98.860 66.205 ;
        RECT 99.030 65.385 99.260 66.375 ;
        RECT 98.510 65.215 99.260 65.385 ;
        RECT 92.525 64.545 97.870 64.980 ;
        RECT 98.510 64.715 98.765 65.215 ;
        RECT 98.935 64.545 99.265 65.045 ;
        RECT 99.435 64.715 99.605 66.835 ;
        RECT 99.965 66.735 100.295 67.095 ;
        RECT 100.465 66.705 100.960 66.875 ;
        RECT 101.165 66.705 102.020 66.875 ;
        RECT 99.835 65.515 100.295 66.565 ;
        RECT 99.775 64.730 100.100 65.515 ;
        RECT 100.465 65.345 100.635 66.705 ;
        RECT 100.805 65.795 101.155 66.415 ;
        RECT 101.325 66.195 101.680 66.415 ;
        RECT 101.325 65.605 101.495 66.195 ;
        RECT 101.850 65.995 102.020 66.705 ;
        RECT 102.895 66.635 103.225 67.095 ;
        RECT 103.435 66.735 103.785 66.905 ;
        RECT 102.225 66.165 103.015 66.415 ;
        RECT 103.435 66.345 103.695 66.735 ;
        RECT 104.005 66.645 104.955 66.925 ;
        RECT 105.125 66.655 105.315 67.095 ;
        RECT 105.485 66.715 106.555 66.885 ;
        RECT 103.185 65.995 103.355 66.175 ;
        RECT 100.465 65.175 100.860 65.345 ;
        RECT 101.030 65.215 101.495 65.605 ;
        RECT 101.665 65.825 103.355 65.995 ;
        RECT 100.690 65.045 100.860 65.175 ;
        RECT 101.665 65.045 101.835 65.825 ;
        RECT 103.525 65.655 103.695 66.345 ;
        RECT 102.195 65.485 103.695 65.655 ;
        RECT 103.885 65.685 104.095 66.475 ;
        RECT 104.265 65.855 104.615 66.475 ;
        RECT 104.785 65.865 104.955 66.645 ;
        RECT 105.485 66.485 105.655 66.715 ;
        RECT 105.125 66.315 105.655 66.485 ;
        RECT 105.125 66.035 105.345 66.315 ;
        RECT 105.825 66.145 106.065 66.545 ;
        RECT 104.785 65.695 105.190 65.865 ;
        RECT 105.525 65.775 106.065 66.145 ;
        RECT 106.235 66.360 106.555 66.715 ;
        RECT 106.800 66.635 107.105 67.095 ;
        RECT 107.275 66.385 107.525 66.915 ;
        RECT 106.235 66.185 106.560 66.360 ;
        RECT 106.235 65.885 107.150 66.185 ;
        RECT 106.410 65.855 107.150 65.885 ;
        RECT 103.885 65.525 104.560 65.685 ;
        RECT 105.020 65.605 105.190 65.695 ;
        RECT 103.885 65.515 104.850 65.525 ;
        RECT 103.525 65.345 103.695 65.485 ;
        RECT 100.270 64.545 100.520 65.005 ;
        RECT 100.690 64.715 100.940 65.045 ;
        RECT 101.155 64.715 101.835 65.045 ;
        RECT 102.005 65.145 103.080 65.315 ;
        RECT 103.525 65.175 104.085 65.345 ;
        RECT 104.390 65.225 104.850 65.515 ;
        RECT 105.020 65.435 106.240 65.605 ;
        RECT 102.005 64.805 102.175 65.145 ;
        RECT 102.410 64.545 102.740 64.975 ;
        RECT 102.910 64.805 103.080 65.145 ;
        RECT 103.375 64.545 103.745 65.005 ;
        RECT 103.915 64.715 104.085 65.175 ;
        RECT 105.020 65.055 105.190 65.435 ;
        RECT 106.410 65.265 106.580 65.855 ;
        RECT 107.320 65.735 107.525 66.385 ;
        RECT 107.695 66.340 107.945 67.095 ;
        RECT 108.225 66.275 108.435 67.095 ;
        RECT 108.605 66.295 108.935 66.925 ;
        RECT 104.320 64.715 105.190 65.055 ;
        RECT 105.780 65.095 106.580 65.265 ;
        RECT 105.360 64.545 105.610 65.005 ;
        RECT 105.780 64.805 105.950 65.095 ;
        RECT 106.130 64.545 106.460 64.925 ;
        RECT 106.800 64.545 107.105 65.685 ;
        RECT 107.275 64.855 107.525 65.735 ;
        RECT 108.605 65.695 108.855 66.295 ;
        RECT 109.105 66.275 109.335 67.095 ;
        RECT 109.545 66.550 114.890 67.095 ;
        RECT 109.025 65.855 109.355 66.105 ;
        RECT 111.130 65.720 111.470 66.550 ;
        RECT 115.105 66.275 115.335 67.095 ;
        RECT 115.505 66.295 115.835 66.925 ;
        RECT 107.695 64.545 107.945 65.685 ;
        RECT 108.225 64.545 108.435 65.685 ;
        RECT 108.605 64.715 108.935 65.695 ;
        RECT 109.105 64.545 109.335 65.685 ;
        RECT 112.950 64.980 113.300 66.230 ;
        RECT 115.085 65.855 115.415 66.105 ;
        RECT 115.585 65.695 115.835 66.295 ;
        RECT 116.005 66.275 116.215 67.095 ;
        RECT 116.905 66.370 117.195 67.095 ;
        RECT 117.365 66.325 120.875 67.095 ;
        RECT 117.365 65.805 119.015 66.325 ;
        RECT 122.025 66.275 122.235 67.095 ;
        RECT 122.405 66.295 122.735 66.925 ;
        RECT 109.545 64.545 114.890 64.980 ;
        RECT 115.105 64.545 115.335 65.685 ;
        RECT 115.505 64.715 115.835 65.695 ;
        RECT 116.005 64.545 116.215 65.685 ;
        RECT 116.905 64.545 117.195 65.710 ;
        RECT 119.185 65.635 120.875 66.155 ;
        RECT 122.405 65.695 122.655 66.295 ;
        RECT 122.905 66.275 123.135 67.095 ;
        RECT 124.270 66.545 124.525 66.835 ;
        RECT 124.695 66.715 125.025 67.095 ;
        RECT 124.270 66.375 125.020 66.545 ;
        RECT 122.825 65.855 123.155 66.105 ;
        RECT 117.365 64.545 120.875 65.635 ;
        RECT 122.025 64.545 122.235 65.685 ;
        RECT 122.405 64.715 122.735 65.695 ;
        RECT 122.905 64.545 123.135 65.685 ;
        RECT 124.270 65.555 124.620 66.205 ;
        RECT 124.790 65.385 125.020 66.375 ;
        RECT 124.270 65.215 125.020 65.385 ;
        RECT 124.270 64.715 124.525 65.215 ;
        RECT 124.695 64.545 125.025 65.045 ;
        RECT 125.195 64.715 125.365 66.835 ;
        RECT 125.725 66.735 126.055 67.095 ;
        RECT 126.225 66.705 126.720 66.875 ;
        RECT 126.925 66.705 127.780 66.875 ;
        RECT 125.595 65.515 126.055 66.565 ;
        RECT 125.535 64.730 125.860 65.515 ;
        RECT 126.225 65.345 126.395 66.705 ;
        RECT 126.565 65.795 126.915 66.415 ;
        RECT 127.085 66.195 127.440 66.415 ;
        RECT 127.085 65.605 127.255 66.195 ;
        RECT 127.610 65.995 127.780 66.705 ;
        RECT 128.655 66.635 128.985 67.095 ;
        RECT 129.195 66.735 129.545 66.905 ;
        RECT 127.985 66.165 128.775 66.415 ;
        RECT 129.195 66.345 129.455 66.735 ;
        RECT 129.765 66.645 130.715 66.925 ;
        RECT 130.885 66.655 131.075 67.095 ;
        RECT 131.245 66.715 132.315 66.885 ;
        RECT 128.945 65.995 129.115 66.175 ;
        RECT 126.225 65.175 126.620 65.345 ;
        RECT 126.790 65.215 127.255 65.605 ;
        RECT 127.425 65.825 129.115 65.995 ;
        RECT 126.450 65.045 126.620 65.175 ;
        RECT 127.425 65.045 127.595 65.825 ;
        RECT 129.285 65.655 129.455 66.345 ;
        RECT 127.955 65.485 129.455 65.655 ;
        RECT 129.645 65.685 129.855 66.475 ;
        RECT 130.025 65.855 130.375 66.475 ;
        RECT 130.545 65.865 130.715 66.645 ;
        RECT 131.245 66.485 131.415 66.715 ;
        RECT 130.885 66.315 131.415 66.485 ;
        RECT 130.885 66.035 131.105 66.315 ;
        RECT 131.585 66.145 131.825 66.545 ;
        RECT 130.545 65.695 130.950 65.865 ;
        RECT 131.285 65.775 131.825 66.145 ;
        RECT 131.995 66.360 132.315 66.715 ;
        RECT 132.560 66.635 132.865 67.095 ;
        RECT 133.035 66.385 133.290 66.915 ;
        RECT 133.930 66.565 134.220 66.915 ;
        RECT 134.415 66.735 134.745 67.095 ;
        RECT 134.915 66.565 135.145 66.870 ;
        RECT 133.930 66.395 135.145 66.565 ;
        RECT 135.335 66.415 135.505 66.790 ;
        RECT 131.995 66.185 132.320 66.360 ;
        RECT 131.995 65.885 132.910 66.185 ;
        RECT 132.170 65.855 132.910 65.885 ;
        RECT 129.645 65.525 130.320 65.685 ;
        RECT 130.780 65.605 130.950 65.695 ;
        RECT 129.645 65.515 130.610 65.525 ;
        RECT 129.285 65.345 129.455 65.485 ;
        RECT 126.030 64.545 126.280 65.005 ;
        RECT 126.450 64.715 126.700 65.045 ;
        RECT 126.915 64.715 127.595 65.045 ;
        RECT 127.765 65.145 128.840 65.315 ;
        RECT 129.285 65.175 129.845 65.345 ;
        RECT 130.150 65.225 130.610 65.515 ;
        RECT 130.780 65.435 132.000 65.605 ;
        RECT 127.765 64.805 127.935 65.145 ;
        RECT 128.170 64.545 128.500 64.975 ;
        RECT 128.670 64.805 128.840 65.145 ;
        RECT 129.135 64.545 129.505 65.005 ;
        RECT 129.675 64.715 129.845 65.175 ;
        RECT 130.780 65.055 130.950 65.435 ;
        RECT 132.170 65.265 132.340 65.855 ;
        RECT 133.080 65.735 133.290 66.385 ;
        RECT 135.335 66.245 135.535 66.415 ;
        RECT 135.765 66.325 137.435 67.095 ;
        RECT 135.335 66.225 135.505 66.245 ;
        RECT 133.990 66.075 134.250 66.185 ;
        RECT 133.985 65.905 134.250 66.075 ;
        RECT 133.990 65.855 134.250 65.905 ;
        RECT 134.430 65.855 134.815 66.185 ;
        RECT 134.985 66.055 135.505 66.225 ;
        RECT 130.080 64.715 130.950 65.055 ;
        RECT 131.540 65.095 132.340 65.265 ;
        RECT 131.120 64.545 131.370 65.005 ;
        RECT 131.540 64.805 131.710 65.095 ;
        RECT 131.890 64.545 132.220 64.925 ;
        RECT 132.560 64.545 132.865 65.685 ;
        RECT 133.035 64.855 133.290 65.735 ;
        RECT 133.930 64.545 134.250 65.685 ;
        RECT 134.430 64.805 134.625 65.855 ;
        RECT 134.985 65.675 135.155 66.055 ;
        RECT 134.805 65.395 135.155 65.675 ;
        RECT 135.345 65.525 135.590 65.885 ;
        RECT 135.765 65.805 136.515 66.325 ;
        RECT 138.065 66.295 138.405 66.925 ;
        RECT 138.695 66.635 138.865 67.095 ;
        RECT 139.135 66.465 139.465 66.910 ;
        RECT 136.685 65.635 137.435 66.155 ;
        RECT 134.805 64.715 135.135 65.395 ;
        RECT 135.335 64.545 135.590 65.345 ;
        RECT 135.765 64.545 137.435 65.635 ;
        RECT 138.065 65.725 138.335 66.295 ;
        RECT 138.715 66.275 139.465 66.465 ;
        RECT 139.635 66.445 139.805 66.765 ;
        RECT 140.030 66.635 140.360 67.095 ;
        RECT 140.560 66.445 140.890 66.925 ;
        RECT 141.105 66.635 141.435 67.095 ;
        RECT 141.605 66.445 141.935 66.925 ;
        RECT 139.635 66.275 141.935 66.445 ;
        RECT 142.665 66.370 142.955 67.095 ;
        RECT 138.715 66.105 139.085 66.275 ;
        RECT 143.240 66.180 143.410 67.095 ;
        RECT 143.580 66.420 143.855 66.765 ;
        RECT 144.045 66.695 144.425 67.095 ;
        RECT 144.595 66.525 144.765 66.875 ;
        RECT 144.935 66.695 145.265 67.095 ;
        RECT 145.465 66.525 145.635 66.875 ;
        RECT 145.835 66.595 146.170 67.095 ;
        RECT 138.505 65.895 139.085 66.105 ;
        RECT 139.255 65.895 139.675 66.105 ;
        RECT 138.825 65.725 139.085 65.895 ;
        RECT 138.065 64.715 138.590 65.725 ;
        RECT 138.825 65.435 139.575 65.725 ;
        RECT 138.825 64.545 139.155 65.265 ;
        RECT 139.325 64.715 139.575 65.435 ;
        RECT 139.845 64.790 140.175 66.105 ;
        RECT 140.385 64.790 140.715 66.105 ;
        RECT 140.885 64.790 141.255 66.105 ;
        RECT 141.465 65.855 141.975 66.105 ;
        RECT 141.585 64.545 141.915 65.665 ;
        RECT 142.665 64.545 142.955 65.710 ;
        RECT 143.240 64.545 143.410 65.725 ;
        RECT 143.580 65.685 143.750 66.420 ;
        RECT 144.025 66.355 145.635 66.525 ;
        RECT 144.025 66.185 144.195 66.355 ;
        RECT 143.920 65.855 144.195 66.185 ;
        RECT 144.365 65.855 144.770 66.185 ;
        RECT 144.025 65.685 144.195 65.855 ;
        RECT 143.580 64.715 143.855 65.685 ;
        RECT 144.025 65.515 144.750 65.685 ;
        RECT 144.940 65.565 145.650 66.185 ;
        RECT 145.820 65.855 146.175 66.425 ;
        RECT 146.345 66.325 149.855 67.095 ;
        RECT 150.945 66.345 152.155 67.095 ;
        RECT 146.345 65.805 147.995 66.325 ;
        RECT 144.580 65.395 144.750 65.515 ;
        RECT 145.850 65.395 146.175 65.685 ;
        RECT 148.165 65.635 149.855 66.155 ;
        RECT 144.065 64.545 144.345 65.345 ;
        RECT 144.580 65.225 146.175 65.395 ;
        RECT 144.515 64.765 146.175 65.055 ;
        RECT 146.345 64.545 149.855 65.635 ;
        RECT 150.945 65.635 151.465 66.175 ;
        RECT 151.635 65.805 152.155 66.345 ;
        RECT 150.945 64.545 152.155 65.635 ;
        RECT 91.060 64.375 152.240 64.545 ;
        RECT 33.585 64.160 35.445 64.330 ;
        RECT 33.585 63.600 33.755 64.160 ;
        RECT 35.275 62.305 35.445 64.160 ;
        RECT 91.145 63.285 92.355 64.375 ;
        RECT 31.705 62.135 35.445 62.305 ;
        RECT 91.145 62.575 91.665 63.115 ;
        RECT 91.835 62.745 92.355 63.285 ;
        RECT 92.575 63.235 92.825 64.375 ;
        RECT 92.995 63.185 93.245 64.065 ;
        RECT 93.415 63.235 93.720 64.375 ;
        RECT 94.060 63.995 94.390 64.375 ;
        RECT 94.570 63.825 94.740 64.115 ;
        RECT 94.910 63.915 95.160 64.375 ;
        RECT 93.940 63.655 94.740 63.825 ;
        RECT 95.330 63.865 96.200 64.205 ;
        RECT 32.650 61.770 32.930 61.850 ;
        RECT 91.145 61.825 92.355 62.575 ;
        RECT 92.575 61.825 92.825 62.580 ;
        RECT 92.995 62.535 93.200 63.185 ;
        RECT 93.940 63.065 94.110 63.655 ;
        RECT 95.330 63.485 95.500 63.865 ;
        RECT 96.435 63.745 96.605 64.205 ;
        RECT 96.775 63.915 97.145 64.375 ;
        RECT 97.440 63.775 97.610 64.115 ;
        RECT 97.780 63.945 98.110 64.375 ;
        RECT 98.345 63.775 98.515 64.115 ;
        RECT 94.280 63.315 95.500 63.485 ;
        RECT 95.670 63.405 96.130 63.695 ;
        RECT 96.435 63.575 96.995 63.745 ;
        RECT 97.440 63.605 98.515 63.775 ;
        RECT 98.685 63.875 99.365 64.205 ;
        RECT 99.580 63.875 99.830 64.205 ;
        RECT 100.000 63.915 100.250 64.375 ;
        RECT 96.825 63.435 96.995 63.575 ;
        RECT 95.670 63.395 96.635 63.405 ;
        RECT 95.330 63.225 95.500 63.315 ;
        RECT 95.960 63.235 96.635 63.395 ;
        RECT 93.370 63.035 94.110 63.065 ;
        RECT 93.370 62.735 94.285 63.035 ;
        RECT 93.960 62.560 94.285 62.735 ;
        RECT 92.995 62.005 93.245 62.535 ;
        RECT 93.415 61.825 93.720 62.285 ;
        RECT 93.965 62.205 94.285 62.560 ;
        RECT 94.455 62.775 94.995 63.145 ;
        RECT 95.330 63.055 95.735 63.225 ;
        RECT 94.455 62.375 94.695 62.775 ;
        RECT 95.175 62.605 95.395 62.885 ;
        RECT 94.865 62.435 95.395 62.605 ;
        RECT 94.865 62.205 95.035 62.435 ;
        RECT 95.565 62.275 95.735 63.055 ;
        RECT 95.905 62.445 96.255 63.065 ;
        RECT 96.425 62.445 96.635 63.235 ;
        RECT 96.825 63.265 98.325 63.435 ;
        RECT 96.825 62.575 96.995 63.265 ;
        RECT 98.685 63.095 98.855 63.875 ;
        RECT 99.660 63.745 99.830 63.875 ;
        RECT 97.165 62.925 98.855 63.095 ;
        RECT 99.025 63.315 99.490 63.705 ;
        RECT 99.660 63.575 100.055 63.745 ;
        RECT 97.165 62.745 97.335 62.925 ;
        RECT 93.965 62.035 95.035 62.205 ;
        RECT 95.205 61.825 95.395 62.265 ;
        RECT 95.565 61.995 96.515 62.275 ;
        RECT 96.825 62.185 97.085 62.575 ;
        RECT 97.505 62.505 98.295 62.755 ;
        RECT 96.735 62.015 97.085 62.185 ;
        RECT 97.295 61.825 97.625 62.285 ;
        RECT 98.500 62.215 98.670 62.925 ;
        RECT 99.025 62.725 99.195 63.315 ;
        RECT 98.840 62.505 99.195 62.725 ;
        RECT 99.365 62.505 99.715 63.125 ;
        RECT 99.885 62.215 100.055 63.575 ;
        RECT 100.420 63.405 100.745 64.190 ;
        RECT 100.225 62.355 100.685 63.405 ;
        RECT 98.500 62.045 99.355 62.215 ;
        RECT 99.560 62.045 100.055 62.215 ;
        RECT 100.225 61.825 100.555 62.185 ;
        RECT 100.915 62.085 101.085 64.205 ;
        RECT 101.255 63.875 101.585 64.375 ;
        RECT 101.755 63.705 102.010 64.205 ;
        RECT 101.260 63.535 102.010 63.705 ;
        RECT 101.260 62.545 101.490 63.535 ;
        RECT 101.660 62.715 102.010 63.365 ;
        RECT 102.245 63.235 102.455 64.375 ;
        RECT 102.625 63.225 102.955 64.205 ;
        RECT 103.125 63.235 103.355 64.375 ;
        RECT 101.260 62.375 102.010 62.545 ;
        RECT 101.255 61.825 101.585 62.205 ;
        RECT 101.755 62.085 102.010 62.375 ;
        RECT 102.245 61.825 102.455 62.645 ;
        RECT 102.625 62.625 102.875 63.225 ;
        RECT 104.025 63.210 104.315 64.375 ;
        RECT 104.485 63.285 105.695 64.375 ;
        RECT 103.045 62.815 103.375 63.065 ;
        RECT 102.625 61.995 102.955 62.625 ;
        RECT 103.125 61.825 103.355 62.645 ;
        RECT 104.485 62.575 105.005 63.115 ;
        RECT 105.175 62.745 105.695 63.285 ;
        RECT 105.865 63.235 106.125 64.205 ;
        RECT 106.320 63.965 106.650 64.375 ;
        RECT 106.850 63.785 107.020 64.205 ;
        RECT 107.235 63.965 107.905 64.375 ;
        RECT 108.140 63.785 108.310 64.205 ;
        RECT 108.615 63.935 108.945 64.375 ;
        RECT 106.295 63.615 108.310 63.785 ;
        RECT 109.115 63.755 109.290 64.205 ;
        RECT 104.025 61.825 104.315 62.550 ;
        RECT 104.485 61.825 105.695 62.575 ;
        RECT 105.865 62.545 106.035 63.235 ;
        RECT 106.295 63.065 106.465 63.615 ;
        RECT 106.205 62.735 106.465 63.065 ;
        RECT 105.865 62.080 106.205 62.545 ;
        RECT 106.635 62.405 106.975 63.435 ;
        RECT 107.165 62.335 107.435 63.435 ;
        RECT 105.870 62.035 106.205 62.080 ;
        RECT 106.375 61.825 106.705 62.205 ;
        RECT 107.165 62.165 107.475 62.335 ;
        RECT 107.165 62.160 107.435 62.165 ;
        RECT 107.660 62.160 107.940 63.435 ;
        RECT 108.140 62.325 108.310 63.615 ;
        RECT 108.660 63.585 109.290 63.755 ;
        RECT 108.660 63.065 108.830 63.585 ;
        RECT 108.480 62.735 108.830 63.065 ;
        RECT 109.010 62.735 109.375 63.415 ;
        RECT 109.565 63.320 109.870 64.105 ;
        RECT 110.050 63.905 110.735 64.375 ;
        RECT 110.045 63.385 110.740 63.695 ;
        RECT 108.660 62.565 108.830 62.735 ;
        RECT 108.660 62.395 109.290 62.565 ;
        RECT 108.140 61.995 108.370 62.325 ;
        RECT 108.615 61.825 108.945 62.205 ;
        RECT 109.115 61.995 109.290 62.395 ;
        RECT 109.565 62.515 109.740 63.320 ;
        RECT 110.915 63.215 111.200 64.160 ;
        RECT 111.375 63.925 111.705 64.375 ;
        RECT 111.875 63.755 112.045 64.185 ;
        RECT 110.340 63.065 111.200 63.215 ;
        RECT 109.915 63.045 111.200 63.065 ;
        RECT 111.370 63.525 112.045 63.755 ;
        RECT 112.770 63.705 113.025 64.205 ;
        RECT 113.195 63.875 113.525 64.375 ;
        RECT 112.770 63.535 113.520 63.705 ;
        RECT 109.915 62.685 110.900 63.045 ;
        RECT 111.370 62.875 111.605 63.525 ;
        RECT 109.565 61.995 109.805 62.515 ;
        RECT 110.730 62.350 110.900 62.685 ;
        RECT 111.070 62.545 111.605 62.875 ;
        RECT 111.385 62.395 111.605 62.545 ;
        RECT 111.775 62.505 112.075 63.355 ;
        RECT 112.770 62.715 113.120 63.365 ;
        RECT 113.290 62.545 113.520 63.535 ;
        RECT 109.975 61.825 110.370 62.320 ;
        RECT 110.730 62.155 111.105 62.350 ;
        RECT 110.935 62.010 111.105 62.155 ;
        RECT 111.385 62.020 111.625 62.395 ;
        RECT 112.770 62.375 113.520 62.545 ;
        RECT 111.795 61.825 112.130 62.330 ;
        RECT 112.770 62.085 113.025 62.375 ;
        RECT 113.195 61.825 113.525 62.205 ;
        RECT 113.695 62.085 113.865 64.205 ;
        RECT 114.035 63.405 114.360 64.190 ;
        RECT 114.530 63.915 114.780 64.375 ;
        RECT 114.950 63.875 115.200 64.205 ;
        RECT 115.415 63.875 116.095 64.205 ;
        RECT 114.950 63.745 115.120 63.875 ;
        RECT 114.725 63.575 115.120 63.745 ;
        RECT 114.095 62.355 114.555 63.405 ;
        RECT 114.725 62.215 114.895 63.575 ;
        RECT 115.290 63.315 115.755 63.705 ;
        RECT 115.065 62.505 115.415 63.125 ;
        RECT 115.585 62.725 115.755 63.315 ;
        RECT 115.925 63.095 116.095 63.875 ;
        RECT 116.265 63.775 116.435 64.115 ;
        RECT 116.670 63.945 117.000 64.375 ;
        RECT 117.170 63.775 117.340 64.115 ;
        RECT 117.635 63.915 118.005 64.375 ;
        RECT 116.265 63.605 117.340 63.775 ;
        RECT 118.175 63.745 118.345 64.205 ;
        RECT 118.580 63.865 119.450 64.205 ;
        RECT 119.620 63.915 119.870 64.375 ;
        RECT 117.785 63.575 118.345 63.745 ;
        RECT 117.785 63.435 117.955 63.575 ;
        RECT 116.455 63.265 117.955 63.435 ;
        RECT 118.650 63.405 119.110 63.695 ;
        RECT 115.925 62.925 117.615 63.095 ;
        RECT 115.585 62.505 115.940 62.725 ;
        RECT 116.110 62.215 116.280 62.925 ;
        RECT 116.485 62.505 117.275 62.755 ;
        RECT 117.445 62.745 117.615 62.925 ;
        RECT 117.785 62.575 117.955 63.265 ;
        RECT 114.225 61.825 114.555 62.185 ;
        RECT 114.725 62.045 115.220 62.215 ;
        RECT 115.425 62.045 116.280 62.215 ;
        RECT 117.155 61.825 117.485 62.285 ;
        RECT 117.695 62.185 117.955 62.575 ;
        RECT 118.145 63.395 119.110 63.405 ;
        RECT 119.280 63.485 119.450 63.865 ;
        RECT 120.040 63.825 120.210 64.115 ;
        RECT 120.390 63.995 120.720 64.375 ;
        RECT 120.040 63.655 120.840 63.825 ;
        RECT 118.145 63.235 118.820 63.395 ;
        RECT 119.280 63.315 120.500 63.485 ;
        RECT 118.145 62.445 118.355 63.235 ;
        RECT 119.280 63.225 119.450 63.315 ;
        RECT 118.525 62.445 118.875 63.065 ;
        RECT 119.045 63.055 119.450 63.225 ;
        RECT 119.045 62.275 119.215 63.055 ;
        RECT 119.385 62.605 119.605 62.885 ;
        RECT 119.785 62.775 120.325 63.145 ;
        RECT 120.670 63.065 120.840 63.655 ;
        RECT 121.060 63.235 121.365 64.375 ;
        RECT 121.535 63.185 121.790 64.065 ;
        RECT 120.670 63.035 121.410 63.065 ;
        RECT 119.385 62.435 119.915 62.605 ;
        RECT 117.695 62.015 118.045 62.185 ;
        RECT 118.265 61.995 119.215 62.275 ;
        RECT 119.385 61.825 119.575 62.265 ;
        RECT 119.745 62.205 119.915 62.435 ;
        RECT 120.085 62.375 120.325 62.775 ;
        RECT 120.495 62.735 121.410 63.035 ;
        RECT 120.495 62.560 120.820 62.735 ;
        RECT 120.495 62.205 120.815 62.560 ;
        RECT 121.580 62.535 121.790 63.185 ;
        RECT 119.745 62.035 120.815 62.205 ;
        RECT 121.060 61.825 121.365 62.285 ;
        RECT 121.535 62.005 121.790 62.535 ;
        RECT 121.965 63.235 122.350 64.205 ;
        RECT 122.520 63.915 122.845 64.375 ;
        RECT 123.365 63.745 123.645 64.205 ;
        RECT 122.520 63.525 123.645 63.745 ;
        RECT 121.965 62.565 122.245 63.235 ;
        RECT 122.520 63.065 122.970 63.525 ;
        RECT 123.835 63.355 124.235 64.205 ;
        RECT 124.635 63.915 124.905 64.375 ;
        RECT 125.075 63.745 125.360 64.205 ;
        RECT 122.415 62.735 122.970 63.065 ;
        RECT 123.140 62.795 124.235 63.355 ;
        RECT 122.520 62.625 122.970 62.735 ;
        RECT 121.965 61.995 122.350 62.565 ;
        RECT 122.520 62.455 123.645 62.625 ;
        RECT 122.520 61.825 122.845 62.285 ;
        RECT 123.365 61.995 123.645 62.455 ;
        RECT 123.835 61.995 124.235 62.795 ;
        RECT 124.405 63.525 125.360 63.745 ;
        RECT 124.405 62.625 124.615 63.525 ;
        RECT 124.785 62.795 125.475 63.355 ;
        RECT 126.605 63.235 126.835 64.375 ;
        RECT 127.005 63.225 127.335 64.205 ;
        RECT 127.505 63.235 127.715 64.375 ;
        RECT 127.945 63.285 129.615 64.375 ;
        RECT 126.585 62.815 126.915 63.065 ;
        RECT 124.405 62.455 125.360 62.625 ;
        RECT 124.635 61.825 124.905 62.285 ;
        RECT 125.075 61.995 125.360 62.455 ;
        RECT 126.605 61.825 126.835 62.645 ;
        RECT 127.085 62.625 127.335 63.225 ;
        RECT 127.005 61.995 127.335 62.625 ;
        RECT 127.505 61.825 127.715 62.645 ;
        RECT 127.945 62.595 128.695 63.115 ;
        RECT 128.865 62.765 129.615 63.285 ;
        RECT 129.785 63.210 130.075 64.375 ;
        RECT 130.245 63.940 135.590 64.375 ;
        RECT 135.765 63.940 141.110 64.375 ;
        RECT 127.945 61.825 129.615 62.595 ;
        RECT 129.785 61.825 130.075 62.550 ;
        RECT 131.830 62.370 132.170 63.200 ;
        RECT 133.650 62.690 134.000 63.940 ;
        RECT 137.350 62.370 137.690 63.200 ;
        RECT 139.170 62.690 139.520 63.940 ;
        RECT 142.215 63.405 142.545 64.190 ;
        RECT 142.215 63.235 142.895 63.405 ;
        RECT 143.075 63.235 143.405 64.375 ;
        RECT 143.585 63.285 146.175 64.375 ;
        RECT 142.205 62.815 142.555 63.065 ;
        RECT 142.725 62.635 142.895 63.235 ;
        RECT 143.065 62.815 143.415 63.065 ;
        RECT 130.245 61.825 135.590 62.370 ;
        RECT 135.765 61.825 141.110 62.370 ;
        RECT 142.225 61.825 142.465 62.635 ;
        RECT 142.635 61.995 142.965 62.635 ;
        RECT 143.135 61.825 143.405 62.635 ;
        RECT 143.585 62.595 144.795 63.115 ;
        RECT 144.965 62.765 146.175 63.285 ;
        RECT 146.405 63.235 146.615 64.375 ;
        RECT 146.785 63.225 147.115 64.205 ;
        RECT 147.285 63.235 147.515 64.375 ;
        RECT 147.725 63.285 150.315 64.375 ;
        RECT 143.585 61.825 146.175 62.595 ;
        RECT 146.405 61.825 146.615 62.645 ;
        RECT 146.785 62.625 147.035 63.225 ;
        RECT 147.205 62.815 147.535 63.065 ;
        RECT 146.785 61.995 147.115 62.625 ;
        RECT 147.285 61.825 147.515 62.645 ;
        RECT 147.725 62.595 148.935 63.115 ;
        RECT 149.105 62.765 150.315 63.285 ;
        RECT 150.945 63.285 152.155 64.375 ;
        RECT 150.945 62.745 151.465 63.285 ;
        RECT 147.725 61.825 150.315 62.595 ;
        RECT 151.635 62.575 152.155 63.115 ;
        RECT 150.945 61.825 152.155 62.575 ;
        RECT 30.400 61.600 32.930 61.770 ;
        RECT 91.060 61.655 152.240 61.825 ;
        RECT 32.650 61.535 32.930 61.600 ;
        RECT 91.145 60.905 92.355 61.655 ;
        RECT 91.145 60.365 91.665 60.905 ;
        RECT 92.525 60.885 96.035 61.655 ;
        RECT 91.835 60.195 92.355 60.735 ;
        RECT 92.525 60.365 94.175 60.885 ;
        RECT 97.125 60.855 97.435 61.655 ;
        RECT 97.640 60.855 98.335 61.485 ;
        RECT 98.710 60.875 99.210 61.485 ;
        RECT 97.640 60.805 97.815 60.855 ;
        RECT 94.345 60.195 96.035 60.715 ;
        RECT 97.135 60.415 97.470 60.685 ;
        RECT 97.640 60.255 97.810 60.805 ;
        RECT 97.980 60.415 98.315 60.665 ;
        RECT 98.505 60.415 98.855 60.665 ;
        RECT 29.750 59.205 30.145 59.570 ;
        RECT 91.145 59.105 92.355 60.195 ;
        RECT 92.525 59.105 96.035 60.195 ;
        RECT 97.125 59.105 97.405 60.245 ;
        RECT 97.575 59.275 97.905 60.255 ;
        RECT 99.040 60.245 99.210 60.875 ;
        RECT 99.840 61.005 100.170 61.485 ;
        RECT 100.340 61.195 100.565 61.655 ;
        RECT 100.735 61.005 101.065 61.485 ;
        RECT 99.840 60.835 101.065 61.005 ;
        RECT 101.255 60.855 101.505 61.655 ;
        RECT 101.675 60.855 102.015 61.485 ;
        RECT 99.380 60.465 99.710 60.665 ;
        RECT 99.880 60.465 100.210 60.665 ;
        RECT 100.380 60.465 100.800 60.665 ;
        RECT 100.975 60.495 101.670 60.665 ;
        RECT 100.975 60.245 101.145 60.495 ;
        RECT 101.840 60.245 102.015 60.855 ;
        RECT 98.075 59.105 98.335 60.245 ;
        RECT 98.710 60.075 101.145 60.245 ;
        RECT 98.710 59.275 99.040 60.075 ;
        RECT 99.210 59.105 99.540 59.905 ;
        RECT 99.840 59.275 100.170 60.075 ;
        RECT 100.815 59.105 101.065 59.905 ;
        RECT 101.335 59.105 101.505 60.245 ;
        RECT 101.675 59.275 102.015 60.245 ;
        RECT 102.185 61.005 102.445 61.485 ;
        RECT 102.615 61.195 102.945 61.655 ;
        RECT 103.135 61.015 103.335 61.435 ;
        RECT 102.185 59.975 102.355 61.005 ;
        RECT 102.525 60.315 102.755 60.745 ;
        RECT 102.925 60.495 103.335 61.015 ;
        RECT 103.505 61.170 104.295 61.435 ;
        RECT 103.505 60.315 103.760 61.170 ;
        RECT 104.475 60.835 104.805 61.255 ;
        RECT 104.975 60.835 105.235 61.655 ;
        RECT 104.475 60.745 104.725 60.835 ;
        RECT 103.930 60.495 104.725 60.745 ;
        RECT 102.525 60.145 104.315 60.315 ;
        RECT 102.185 59.275 102.460 59.975 ;
        RECT 102.630 59.850 103.345 60.145 ;
        RECT 103.565 59.785 103.895 59.975 ;
        RECT 102.670 59.105 102.885 59.650 ;
        RECT 103.055 59.275 103.530 59.615 ;
        RECT 103.700 59.610 103.895 59.785 ;
        RECT 104.065 59.780 104.315 60.145 ;
        RECT 103.700 59.105 104.315 59.610 ;
        RECT 104.555 59.275 104.725 60.495 ;
        RECT 104.895 59.785 105.235 60.665 ;
        RECT 104.975 59.105 105.235 59.615 ;
        RECT 105.415 59.285 105.675 61.475 ;
        RECT 105.935 61.285 106.605 61.655 ;
        RECT 106.785 61.105 107.095 61.475 ;
        RECT 105.865 60.905 107.095 61.105 ;
        RECT 105.865 60.235 106.155 60.905 ;
        RECT 107.275 60.725 107.505 61.365 ;
        RECT 107.685 60.925 107.975 61.655 ;
        RECT 108.165 61.110 113.510 61.655 ;
        RECT 106.335 60.415 106.800 60.725 ;
        RECT 106.980 60.415 107.505 60.725 ;
        RECT 107.685 60.415 107.985 60.745 ;
        RECT 109.750 60.280 110.090 61.110 ;
        RECT 105.865 60.015 106.635 60.235 ;
        RECT 105.845 59.105 106.185 59.835 ;
        RECT 106.365 59.285 106.635 60.015 ;
        RECT 106.815 59.995 107.975 60.235 ;
        RECT 106.815 59.285 107.045 59.995 ;
        RECT 107.215 59.105 107.545 59.815 ;
        RECT 107.715 59.285 107.975 59.995 ;
        RECT 111.570 59.540 111.920 60.790 ;
        RECT 108.165 59.105 113.510 59.540 ;
        RECT 114.155 59.285 114.415 61.475 ;
        RECT 114.675 61.285 115.345 61.655 ;
        RECT 115.525 61.105 115.835 61.475 ;
        RECT 114.605 60.905 115.835 61.105 ;
        RECT 114.605 60.235 114.895 60.905 ;
        RECT 116.015 60.725 116.245 61.365 ;
        RECT 116.425 60.925 116.715 61.655 ;
        RECT 116.905 60.930 117.195 61.655 ;
        RECT 117.365 61.145 117.670 61.655 ;
        RECT 115.075 60.415 115.540 60.725 ;
        RECT 115.720 60.415 116.245 60.725 ;
        RECT 116.425 60.415 116.725 60.745 ;
        RECT 117.365 60.415 117.680 60.975 ;
        RECT 117.850 60.665 118.100 61.475 ;
        RECT 118.270 61.130 118.530 61.655 ;
        RECT 118.710 60.665 118.960 61.475 ;
        RECT 119.130 61.095 119.390 61.655 ;
        RECT 119.560 61.005 119.820 61.460 ;
        RECT 119.990 61.175 120.250 61.655 ;
        RECT 120.420 61.005 120.680 61.460 ;
        RECT 120.850 61.175 121.110 61.655 ;
        RECT 121.280 61.005 121.540 61.460 ;
        RECT 121.710 61.175 121.955 61.655 ;
        RECT 122.125 61.005 122.400 61.460 ;
        RECT 122.570 61.175 122.815 61.655 ;
        RECT 122.985 61.005 123.245 61.460 ;
        RECT 123.425 61.175 123.675 61.655 ;
        RECT 123.845 61.005 124.105 61.460 ;
        RECT 124.285 61.175 124.535 61.655 ;
        RECT 124.705 61.005 124.965 61.460 ;
        RECT 125.145 61.175 125.405 61.655 ;
        RECT 125.575 61.005 125.835 61.460 ;
        RECT 126.005 61.175 126.305 61.655 ;
        RECT 126.565 61.110 131.910 61.655 ;
        RECT 132.085 61.110 137.430 61.655 ;
        RECT 119.560 60.835 126.305 61.005 ;
        RECT 117.850 60.415 124.970 60.665 ;
        RECT 114.605 60.015 115.375 60.235 ;
        RECT 114.585 59.105 114.925 59.835 ;
        RECT 115.105 59.285 115.375 60.015 ;
        RECT 115.555 59.995 116.715 60.235 ;
        RECT 115.555 59.285 115.785 59.995 ;
        RECT 115.955 59.105 116.285 59.815 ;
        RECT 116.455 59.285 116.715 59.995 ;
        RECT 116.905 59.105 117.195 60.270 ;
        RECT 117.375 59.105 117.670 59.915 ;
        RECT 117.850 59.275 118.095 60.415 ;
        RECT 118.270 59.105 118.530 59.915 ;
        RECT 118.710 59.280 118.960 60.415 ;
        RECT 125.140 60.245 126.305 60.835 ;
        RECT 128.150 60.280 128.490 61.110 ;
        RECT 119.560 60.020 126.305 60.245 ;
        RECT 119.560 60.005 124.965 60.020 ;
        RECT 119.130 59.110 119.390 59.905 ;
        RECT 119.560 59.280 119.820 60.005 ;
        RECT 119.990 59.110 120.250 59.835 ;
        RECT 120.420 59.280 120.680 60.005 ;
        RECT 120.850 59.110 121.110 59.835 ;
        RECT 121.280 59.280 121.540 60.005 ;
        RECT 121.710 59.110 121.970 59.835 ;
        RECT 122.140 59.280 122.400 60.005 ;
        RECT 122.570 59.110 122.815 59.835 ;
        RECT 122.985 59.280 123.245 60.005 ;
        RECT 123.430 59.110 123.675 59.835 ;
        RECT 123.845 59.280 124.105 60.005 ;
        RECT 124.290 59.110 124.535 59.835 ;
        RECT 124.705 59.280 124.965 60.005 ;
        RECT 125.150 59.110 125.405 59.835 ;
        RECT 125.575 59.280 125.865 60.020 ;
        RECT 119.130 59.105 125.405 59.110 ;
        RECT 126.035 59.105 126.305 59.850 ;
        RECT 129.970 59.540 130.320 60.790 ;
        RECT 133.670 60.280 134.010 61.110 ;
        RECT 137.605 60.885 141.115 61.655 ;
        RECT 141.285 60.905 142.495 61.655 ;
        RECT 142.665 60.930 142.955 61.655 ;
        RECT 135.490 59.540 135.840 60.790 ;
        RECT 137.605 60.365 139.255 60.885 ;
        RECT 139.425 60.195 141.115 60.715 ;
        RECT 141.285 60.365 141.805 60.905 ;
        RECT 143.125 60.885 145.715 61.655 ;
        RECT 141.975 60.195 142.495 60.735 ;
        RECT 143.125 60.365 144.335 60.885 ;
        RECT 145.925 60.835 146.155 61.655 ;
        RECT 146.325 60.855 146.655 61.485 ;
        RECT 126.565 59.105 131.910 59.540 ;
        RECT 132.085 59.105 137.430 59.540 ;
        RECT 137.605 59.105 141.115 60.195 ;
        RECT 141.285 59.105 142.495 60.195 ;
        RECT 142.665 59.105 142.955 60.270 ;
        RECT 144.505 60.195 145.715 60.715 ;
        RECT 145.905 60.415 146.235 60.665 ;
        RECT 146.405 60.255 146.655 60.855 ;
        RECT 146.825 60.835 147.035 61.655 ;
        RECT 147.265 60.915 147.650 61.485 ;
        RECT 147.820 61.195 148.145 61.655 ;
        RECT 148.665 61.025 148.945 61.485 ;
        RECT 143.125 59.105 145.715 60.195 ;
        RECT 145.925 59.105 146.155 60.245 ;
        RECT 146.325 59.275 146.655 60.255 ;
        RECT 147.265 60.245 147.545 60.915 ;
        RECT 147.820 60.855 148.945 61.025 ;
        RECT 147.820 60.745 148.270 60.855 ;
        RECT 147.715 60.415 148.270 60.745 ;
        RECT 149.135 60.685 149.535 61.485 ;
        RECT 149.935 61.195 150.205 61.655 ;
        RECT 150.375 61.025 150.660 61.485 ;
        RECT 146.825 59.105 147.035 60.245 ;
        RECT 147.265 59.275 147.650 60.245 ;
        RECT 147.820 59.955 148.270 60.415 ;
        RECT 148.440 60.125 149.535 60.685 ;
        RECT 147.820 59.735 148.945 59.955 ;
        RECT 147.820 59.105 148.145 59.565 ;
        RECT 148.665 59.275 148.945 59.735 ;
        RECT 149.135 59.275 149.535 60.125 ;
        RECT 149.705 60.855 150.660 61.025 ;
        RECT 150.945 60.905 152.155 61.655 ;
        RECT 149.705 59.955 149.915 60.855 ;
        RECT 150.085 60.125 150.775 60.685 ;
        RECT 150.945 60.195 151.465 60.735 ;
        RECT 151.635 60.365 152.155 60.905 ;
        RECT 149.705 59.735 150.660 59.955 ;
        RECT 149.935 59.105 150.205 59.565 ;
        RECT 150.375 59.275 150.660 59.735 ;
        RECT 150.945 59.105 152.155 60.195 ;
        RECT 28.690 59.090 29.305 59.095 ;
        RECT 91.060 58.935 152.240 59.105 ;
        RECT 26.380 58.165 27.105 58.735 ;
        RECT 25.950 57.995 27.105 58.165 ;
        RECT 26.380 57.705 27.105 57.995 ;
        RECT 91.145 57.845 92.355 58.935 ;
        RECT 92.525 57.845 96.035 58.935 ;
        RECT 96.670 58.135 96.925 58.935 ;
        RECT 97.125 58.085 97.455 58.765 ;
        RECT 6.030 56.670 6.380 57.510 ;
        RECT 7.425 57.345 8.225 57.510 ;
        RECT 22.730 56.360 23.980 57.440 ;
        RECT 91.145 57.135 91.665 57.675 ;
        RECT 91.835 57.305 92.355 57.845 ;
        RECT 92.525 57.155 94.175 57.675 ;
        RECT 94.345 57.325 96.035 57.845 ;
        RECT 96.670 57.595 96.915 57.955 ;
        RECT 97.105 57.805 97.455 58.085 ;
        RECT 97.105 57.425 97.275 57.805 ;
        RECT 97.635 57.625 97.830 58.675 ;
        RECT 98.010 57.795 98.330 58.935 ;
        RECT 98.505 58.215 98.965 58.765 ;
        RECT 99.155 58.215 99.485 58.935 ;
        RECT 96.755 57.255 97.275 57.425 ;
        RECT 97.445 57.295 97.830 57.625 ;
        RECT 98.010 57.575 98.270 57.625 ;
        RECT 98.010 57.405 98.275 57.575 ;
        RECT 98.010 57.295 98.270 57.405 ;
        RECT 91.145 56.385 92.355 57.135 ;
        RECT 92.525 56.385 96.035 57.155 ;
        RECT 96.755 56.895 96.925 57.255 ;
        RECT 96.725 56.725 96.925 56.895 ;
        RECT 96.755 56.690 96.925 56.725 ;
        RECT 97.115 56.915 98.330 57.085 ;
        RECT 97.115 56.610 97.345 56.915 ;
        RECT 97.515 56.385 97.845 56.745 ;
        RECT 98.040 56.565 98.330 56.915 ;
        RECT 98.505 56.845 98.755 58.215 ;
        RECT 99.685 58.045 99.985 58.595 ;
        RECT 100.155 58.265 100.435 58.935 ;
        RECT 99.045 57.875 99.985 58.045 ;
        RECT 100.805 58.215 101.265 58.765 ;
        RECT 101.455 58.215 101.785 58.935 ;
        RECT 99.045 57.625 99.215 57.875 ;
        RECT 100.355 57.625 100.620 57.985 ;
        RECT 98.925 57.295 99.215 57.625 ;
        RECT 99.385 57.375 99.725 57.625 ;
        RECT 99.945 57.375 100.620 57.625 ;
        RECT 99.045 57.205 99.215 57.295 ;
        RECT 99.045 57.015 100.435 57.205 ;
        RECT 98.505 56.555 99.065 56.845 ;
        RECT 99.235 56.385 99.485 56.845 ;
        RECT 100.105 56.655 100.435 57.015 ;
        RECT 100.805 56.845 101.055 58.215 ;
        RECT 101.985 58.045 102.285 58.595 ;
        RECT 102.455 58.265 102.735 58.935 ;
        RECT 101.345 57.875 102.285 58.045 ;
        RECT 101.345 57.625 101.515 57.875 ;
        RECT 102.655 57.625 102.920 57.985 ;
        RECT 104.025 57.770 104.315 58.935 ;
        RECT 104.485 58.500 109.830 58.935 ;
        RECT 101.225 57.295 101.515 57.625 ;
        RECT 101.685 57.375 102.025 57.625 ;
        RECT 102.245 57.375 102.920 57.625 ;
        RECT 101.345 57.205 101.515 57.295 ;
        RECT 101.345 57.015 102.735 57.205 ;
        RECT 100.805 56.555 101.365 56.845 ;
        RECT 101.535 56.385 101.785 56.845 ;
        RECT 102.405 56.655 102.735 57.015 ;
        RECT 104.025 56.385 104.315 57.110 ;
        RECT 106.070 56.930 106.410 57.760 ;
        RECT 107.890 57.250 108.240 58.500 ;
        RECT 110.005 57.845 111.675 58.935 ;
        RECT 111.935 58.190 112.205 58.935 ;
        RECT 112.835 58.930 119.110 58.935 ;
        RECT 112.375 58.020 112.665 58.760 ;
        RECT 112.835 58.205 113.090 58.930 ;
        RECT 113.275 58.035 113.535 58.760 ;
        RECT 113.705 58.205 113.950 58.930 ;
        RECT 114.135 58.035 114.395 58.760 ;
        RECT 114.565 58.205 114.810 58.930 ;
        RECT 114.995 58.035 115.255 58.760 ;
        RECT 115.425 58.205 115.670 58.930 ;
        RECT 115.840 58.035 116.100 58.760 ;
        RECT 116.270 58.205 116.530 58.930 ;
        RECT 116.700 58.035 116.960 58.760 ;
        RECT 117.130 58.205 117.390 58.930 ;
        RECT 117.560 58.035 117.820 58.760 ;
        RECT 117.990 58.205 118.250 58.930 ;
        RECT 118.420 58.035 118.680 58.760 ;
        RECT 118.850 58.135 119.110 58.930 ;
        RECT 113.275 58.020 118.680 58.035 ;
        RECT 110.005 57.155 110.755 57.675 ;
        RECT 110.925 57.325 111.675 57.845 ;
        RECT 111.935 57.795 118.680 58.020 ;
        RECT 111.935 57.205 113.100 57.795 ;
        RECT 119.280 57.625 119.530 58.760 ;
        RECT 119.710 58.125 119.970 58.935 ;
        RECT 120.145 57.625 120.390 58.765 ;
        RECT 120.570 58.125 120.865 58.935 ;
        RECT 121.045 57.845 124.555 58.935 ;
        RECT 113.270 57.375 120.390 57.625 ;
        RECT 104.485 56.385 109.830 56.930 ;
        RECT 110.005 56.385 111.675 57.155 ;
        RECT 111.935 57.035 118.680 57.205 ;
        RECT 111.935 56.385 112.235 56.865 ;
        RECT 112.405 56.580 112.665 57.035 ;
        RECT 112.835 56.385 113.095 56.865 ;
        RECT 113.275 56.580 113.535 57.035 ;
        RECT 113.705 56.385 113.955 56.865 ;
        RECT 114.135 56.580 114.395 57.035 ;
        RECT 114.565 56.385 114.815 56.865 ;
        RECT 114.995 56.580 115.255 57.035 ;
        RECT 115.425 56.385 115.670 56.865 ;
        RECT 115.840 56.580 116.115 57.035 ;
        RECT 116.285 56.385 116.530 56.865 ;
        RECT 116.700 56.580 116.960 57.035 ;
        RECT 117.130 56.385 117.390 56.865 ;
        RECT 117.560 56.580 117.820 57.035 ;
        RECT 117.990 56.385 118.250 56.865 ;
        RECT 118.420 56.580 118.680 57.035 ;
        RECT 118.850 56.385 119.110 56.945 ;
        RECT 119.280 56.565 119.530 57.375 ;
        RECT 119.710 56.385 119.970 56.910 ;
        RECT 120.140 56.565 120.390 57.375 ;
        RECT 120.560 57.065 120.875 57.625 ;
        RECT 121.045 57.155 122.695 57.675 ;
        RECT 122.865 57.325 124.555 57.845 ;
        RECT 125.245 57.795 125.455 58.935 ;
        RECT 125.625 57.785 125.955 58.765 ;
        RECT 126.125 57.795 126.355 58.935 ;
        RECT 126.655 58.005 126.825 58.765 ;
        RECT 127.005 58.175 127.335 58.935 ;
        RECT 126.655 57.835 127.320 58.005 ;
        RECT 127.505 57.860 127.775 58.765 ;
        RECT 120.570 56.385 120.875 56.895 ;
        RECT 121.045 56.385 124.555 57.155 ;
        RECT 125.245 56.385 125.455 57.205 ;
        RECT 125.625 57.185 125.875 57.785 ;
        RECT 127.150 57.690 127.320 57.835 ;
        RECT 126.045 57.375 126.375 57.625 ;
        RECT 126.585 57.285 126.915 57.655 ;
        RECT 127.150 57.360 127.435 57.690 ;
        RECT 125.625 56.555 125.955 57.185 ;
        RECT 126.125 56.385 126.355 57.205 ;
        RECT 127.150 57.105 127.320 57.360 ;
        RECT 126.655 56.935 127.320 57.105 ;
        RECT 127.605 57.060 127.775 57.860 ;
        RECT 127.945 57.845 129.615 58.935 ;
        RECT 126.655 56.555 126.825 56.935 ;
        RECT 127.005 56.385 127.335 56.765 ;
        RECT 127.515 56.555 127.775 57.060 ;
        RECT 127.945 57.155 128.695 57.675 ;
        RECT 128.865 57.325 129.615 57.845 ;
        RECT 129.785 57.770 130.075 58.935 ;
        RECT 130.430 57.965 130.820 58.140 ;
        RECT 131.305 58.135 131.635 58.935 ;
        RECT 131.805 58.145 132.340 58.765 ;
        RECT 130.430 57.795 131.855 57.965 ;
        RECT 127.945 56.385 129.615 57.155 ;
        RECT 129.785 56.385 130.075 57.110 ;
        RECT 130.305 57.065 130.660 57.625 ;
        RECT 130.830 56.895 131.000 57.795 ;
        RECT 131.170 57.065 131.435 57.625 ;
        RECT 131.685 57.295 131.855 57.795 ;
        RECT 132.025 57.125 132.340 58.145 ;
        RECT 130.410 56.385 130.650 56.895 ;
        RECT 130.830 56.565 131.110 56.895 ;
        RECT 131.340 56.385 131.555 56.895 ;
        RECT 131.725 56.555 132.340 57.125 ;
        RECT 133.005 57.860 133.275 58.765 ;
        RECT 133.445 58.175 133.775 58.935 ;
        RECT 133.955 58.005 134.125 58.765 ;
        RECT 134.385 58.500 139.730 58.935 ;
        RECT 133.005 57.060 133.175 57.860 ;
        RECT 133.460 57.835 134.125 58.005 ;
        RECT 133.460 57.690 133.630 57.835 ;
        RECT 133.345 57.360 133.630 57.690 ;
        RECT 133.460 57.105 133.630 57.360 ;
        RECT 133.865 57.285 134.195 57.655 ;
        RECT 133.005 56.555 133.265 57.060 ;
        RECT 133.460 56.935 134.125 57.105 ;
        RECT 133.445 56.385 133.775 56.765 ;
        RECT 133.955 56.555 134.125 56.935 ;
        RECT 135.970 56.930 136.310 57.760 ;
        RECT 137.790 57.250 138.140 58.500 ;
        RECT 139.905 57.845 141.115 58.935 ;
        RECT 141.290 58.265 141.545 58.765 ;
        RECT 141.715 58.435 142.045 58.935 ;
        RECT 141.290 58.095 142.040 58.265 ;
        RECT 139.905 57.135 140.425 57.675 ;
        RECT 140.595 57.305 141.115 57.845 ;
        RECT 141.290 57.275 141.640 57.925 ;
        RECT 134.385 56.385 139.730 56.930 ;
        RECT 139.905 56.385 141.115 57.135 ;
        RECT 141.810 57.105 142.040 58.095 ;
        RECT 141.290 56.935 142.040 57.105 ;
        RECT 141.290 56.645 141.545 56.935 ;
        RECT 141.715 56.385 142.045 56.765 ;
        RECT 142.215 56.645 142.385 58.765 ;
        RECT 142.555 57.965 142.880 58.750 ;
        RECT 143.050 58.475 143.300 58.935 ;
        RECT 143.470 58.435 143.720 58.765 ;
        RECT 143.935 58.435 144.615 58.765 ;
        RECT 143.470 58.305 143.640 58.435 ;
        RECT 143.245 58.135 143.640 58.305 ;
        RECT 142.615 56.915 143.075 57.965 ;
        RECT 143.245 56.775 143.415 58.135 ;
        RECT 143.810 57.875 144.275 58.265 ;
        RECT 143.585 57.065 143.935 57.685 ;
        RECT 144.105 57.285 144.275 57.875 ;
        RECT 144.445 57.655 144.615 58.435 ;
        RECT 144.785 58.335 144.955 58.675 ;
        RECT 145.190 58.505 145.520 58.935 ;
        RECT 145.690 58.335 145.860 58.675 ;
        RECT 146.155 58.475 146.525 58.935 ;
        RECT 144.785 58.165 145.860 58.335 ;
        RECT 146.695 58.305 146.865 58.765 ;
        RECT 147.100 58.425 147.970 58.765 ;
        RECT 148.140 58.475 148.390 58.935 ;
        RECT 146.305 58.135 146.865 58.305 ;
        RECT 146.305 57.995 146.475 58.135 ;
        RECT 144.975 57.825 146.475 57.995 ;
        RECT 147.170 57.965 147.630 58.255 ;
        RECT 144.445 57.485 146.135 57.655 ;
        RECT 144.105 57.065 144.460 57.285 ;
        RECT 144.630 56.775 144.800 57.485 ;
        RECT 145.005 57.065 145.795 57.315 ;
        RECT 145.965 57.305 146.135 57.485 ;
        RECT 146.305 57.135 146.475 57.825 ;
        RECT 142.745 56.385 143.075 56.745 ;
        RECT 143.245 56.605 143.740 56.775 ;
        RECT 143.945 56.605 144.800 56.775 ;
        RECT 145.675 56.385 146.005 56.845 ;
        RECT 146.215 56.745 146.475 57.135 ;
        RECT 146.665 57.955 147.630 57.965 ;
        RECT 147.800 58.045 147.970 58.425 ;
        RECT 148.560 58.385 148.730 58.675 ;
        RECT 148.910 58.555 149.240 58.935 ;
        RECT 148.560 58.215 149.360 58.385 ;
        RECT 146.665 57.795 147.340 57.955 ;
        RECT 147.800 57.875 149.020 58.045 ;
        RECT 146.665 57.005 146.875 57.795 ;
        RECT 147.800 57.785 147.970 57.875 ;
        RECT 147.045 57.005 147.395 57.625 ;
        RECT 147.565 57.615 147.970 57.785 ;
        RECT 147.565 56.835 147.735 57.615 ;
        RECT 147.905 57.165 148.125 57.445 ;
        RECT 148.305 57.335 148.845 57.705 ;
        RECT 149.190 57.625 149.360 58.215 ;
        RECT 149.580 57.795 149.885 58.935 ;
        RECT 150.055 57.745 150.310 58.625 ;
        RECT 149.190 57.595 149.930 57.625 ;
        RECT 147.905 56.995 148.435 57.165 ;
        RECT 146.215 56.575 146.565 56.745 ;
        RECT 146.785 56.555 147.735 56.835 ;
        RECT 147.905 56.385 148.095 56.825 ;
        RECT 148.265 56.765 148.435 56.995 ;
        RECT 148.605 56.935 148.845 57.335 ;
        RECT 149.015 57.295 149.930 57.595 ;
        RECT 149.015 57.120 149.340 57.295 ;
        RECT 149.015 56.765 149.335 57.120 ;
        RECT 150.100 57.095 150.310 57.745 ;
        RECT 150.945 57.845 152.155 58.935 ;
        RECT 150.945 57.305 151.465 57.845 ;
        RECT 151.635 57.135 152.155 57.675 ;
        RECT 148.265 56.595 149.335 56.765 ;
        RECT 149.580 56.385 149.885 56.845 ;
        RECT 150.055 56.565 150.310 57.095 ;
        RECT 150.945 56.385 152.155 57.135 ;
        RECT 91.060 56.215 152.240 56.385 ;
        RECT 6.030 53.590 6.380 55.670 ;
        RECT 91.145 55.465 92.355 56.215 ;
        RECT 92.525 55.670 97.870 56.215 ;
        RECT 91.145 54.925 91.665 55.465 ;
        RECT 91.835 54.755 92.355 55.295 ;
        RECT 94.110 54.840 94.450 55.670 ;
        RECT 98.525 55.405 98.765 56.215 ;
        RECT 98.935 55.405 99.265 56.045 ;
        RECT 99.435 55.405 99.705 56.215 ;
        RECT 99.885 55.670 105.230 56.215 ;
        RECT 105.405 55.670 110.750 56.215 ;
        RECT 91.145 53.665 92.355 54.755 ;
        RECT 95.930 54.100 96.280 55.350 ;
        RECT 98.505 54.975 98.855 55.225 ;
        RECT 99.025 54.805 99.195 55.405 ;
        RECT 99.365 54.975 99.715 55.225 ;
        RECT 101.470 54.840 101.810 55.670 ;
        RECT 98.515 54.635 99.195 54.805 ;
        RECT 92.525 53.665 97.870 54.100 ;
        RECT 98.515 53.850 98.845 54.635 ;
        RECT 99.375 53.665 99.705 54.805 ;
        RECT 103.290 54.100 103.640 55.350 ;
        RECT 106.990 54.840 107.330 55.670 ;
        RECT 110.925 55.465 112.135 56.215 ;
        RECT 108.810 54.100 109.160 55.350 ;
        RECT 110.925 54.925 111.445 55.465 ;
        RECT 112.305 55.395 112.565 56.215 ;
        RECT 112.735 55.395 113.065 55.815 ;
        RECT 113.245 55.730 114.035 55.995 ;
        RECT 112.815 55.305 113.065 55.395 ;
        RECT 111.615 54.755 112.135 55.295 ;
        RECT 99.885 53.665 105.230 54.100 ;
        RECT 105.405 53.665 110.750 54.100 ;
        RECT 110.925 53.665 112.135 54.755 ;
        RECT 112.305 54.345 112.645 55.225 ;
        RECT 112.815 55.055 113.610 55.305 ;
        RECT 112.305 53.665 112.565 54.175 ;
        RECT 112.815 53.835 112.985 55.055 ;
        RECT 113.780 54.875 114.035 55.730 ;
        RECT 114.205 55.575 114.405 55.995 ;
        RECT 114.595 55.755 114.925 56.215 ;
        RECT 114.205 55.055 114.615 55.575 ;
        RECT 115.095 55.565 115.355 56.045 ;
        RECT 114.785 54.875 115.015 55.305 ;
        RECT 113.225 54.705 115.015 54.875 ;
        RECT 113.225 54.340 113.475 54.705 ;
        RECT 113.645 54.345 113.975 54.535 ;
        RECT 114.195 54.410 114.910 54.705 ;
        RECT 115.185 54.535 115.355 55.565 ;
        RECT 113.645 54.170 113.840 54.345 ;
        RECT 113.225 53.665 113.840 54.170 ;
        RECT 114.010 53.835 114.485 54.175 ;
        RECT 114.655 53.665 114.870 54.210 ;
        RECT 115.080 53.835 115.355 54.535 ;
        RECT 115.525 55.540 115.785 56.045 ;
        RECT 115.965 55.835 116.295 56.215 ;
        RECT 116.475 55.665 116.645 56.045 ;
        RECT 115.525 54.740 115.695 55.540 ;
        RECT 115.980 55.495 116.645 55.665 ;
        RECT 115.980 55.240 116.150 55.495 ;
        RECT 116.905 55.490 117.195 56.215 ;
        RECT 118.325 55.395 118.555 56.215 ;
        RECT 118.725 55.415 119.055 56.045 ;
        RECT 115.865 54.910 116.150 55.240 ;
        RECT 116.385 54.945 116.715 55.315 ;
        RECT 118.305 54.975 118.635 55.225 ;
        RECT 115.980 54.765 116.150 54.910 ;
        RECT 115.525 53.835 115.795 54.740 ;
        RECT 115.980 54.595 116.645 54.765 ;
        RECT 115.965 53.665 116.295 54.425 ;
        RECT 116.475 53.835 116.645 54.595 ;
        RECT 116.905 53.665 117.195 54.830 ;
        RECT 118.805 54.815 119.055 55.415 ;
        RECT 119.225 55.395 119.435 56.215 ;
        RECT 119.665 55.445 121.335 56.215 ;
        RECT 121.555 55.460 121.805 56.215 ;
        RECT 121.975 55.505 122.225 56.035 ;
        RECT 122.395 55.755 122.700 56.215 ;
        RECT 122.945 55.835 124.015 56.005 ;
        RECT 119.665 54.925 120.415 55.445 ;
        RECT 118.325 53.665 118.555 54.805 ;
        RECT 118.725 53.835 119.055 54.815 ;
        RECT 119.225 53.665 119.435 54.805 ;
        RECT 120.585 54.755 121.335 55.275 ;
        RECT 121.975 54.855 122.180 55.505 ;
        RECT 122.945 55.480 123.265 55.835 ;
        RECT 122.940 55.305 123.265 55.480 ;
        RECT 122.350 55.005 123.265 55.305 ;
        RECT 123.435 55.265 123.675 55.665 ;
        RECT 123.845 55.605 124.015 55.835 ;
        RECT 124.185 55.775 124.375 56.215 ;
        RECT 124.545 55.765 125.495 56.045 ;
        RECT 125.715 55.855 126.065 56.025 ;
        RECT 123.845 55.435 124.375 55.605 ;
        RECT 122.350 54.975 123.090 55.005 ;
        RECT 119.665 53.665 121.335 54.755 ;
        RECT 121.555 53.665 121.805 54.805 ;
        RECT 121.975 53.975 122.225 54.855 ;
        RECT 122.395 53.665 122.700 54.805 ;
        RECT 122.920 54.385 123.090 54.975 ;
        RECT 123.435 54.895 123.975 55.265 ;
        RECT 124.155 55.155 124.375 55.435 ;
        RECT 124.545 54.985 124.715 55.765 ;
        RECT 124.310 54.815 124.715 54.985 ;
        RECT 124.885 54.975 125.235 55.595 ;
        RECT 124.310 54.725 124.480 54.815 ;
        RECT 125.405 54.805 125.615 55.595 ;
        RECT 123.260 54.555 124.480 54.725 ;
        RECT 124.940 54.645 125.615 54.805 ;
        RECT 122.920 54.215 123.720 54.385 ;
        RECT 123.040 53.665 123.370 54.045 ;
        RECT 123.550 53.925 123.720 54.215 ;
        RECT 124.310 54.175 124.480 54.555 ;
        RECT 124.650 54.635 125.615 54.645 ;
        RECT 125.805 55.465 126.065 55.855 ;
        RECT 126.275 55.755 126.605 56.215 ;
        RECT 127.480 55.825 128.335 55.995 ;
        RECT 128.540 55.825 129.035 55.995 ;
        RECT 129.205 55.855 129.535 56.215 ;
        RECT 125.805 54.775 125.975 55.465 ;
        RECT 126.145 55.115 126.315 55.295 ;
        RECT 126.485 55.285 127.275 55.535 ;
        RECT 127.480 55.115 127.650 55.825 ;
        RECT 127.820 55.315 128.175 55.535 ;
        RECT 126.145 54.945 127.835 55.115 ;
        RECT 124.650 54.345 125.110 54.635 ;
        RECT 125.805 54.605 127.305 54.775 ;
        RECT 125.805 54.465 125.975 54.605 ;
        RECT 125.415 54.295 125.975 54.465 ;
        RECT 123.890 53.665 124.140 54.125 ;
        RECT 124.310 53.835 125.180 54.175 ;
        RECT 125.415 53.835 125.585 54.295 ;
        RECT 126.420 54.265 127.495 54.435 ;
        RECT 125.755 53.665 126.125 54.125 ;
        RECT 126.420 53.925 126.590 54.265 ;
        RECT 126.760 53.665 127.090 54.095 ;
        RECT 127.325 53.925 127.495 54.265 ;
        RECT 127.665 54.165 127.835 54.945 ;
        RECT 128.005 54.725 128.175 55.315 ;
        RECT 128.345 54.915 128.695 55.535 ;
        RECT 128.005 54.335 128.470 54.725 ;
        RECT 128.865 54.465 129.035 55.825 ;
        RECT 129.205 54.635 129.665 55.685 ;
        RECT 128.640 54.295 129.035 54.465 ;
        RECT 128.640 54.165 128.810 54.295 ;
        RECT 127.665 53.835 128.345 54.165 ;
        RECT 128.560 53.835 128.810 54.165 ;
        RECT 128.980 53.665 129.230 54.125 ;
        RECT 129.400 53.850 129.725 54.635 ;
        RECT 129.895 53.835 130.065 55.955 ;
        RECT 130.235 55.835 130.565 56.215 ;
        RECT 130.735 55.665 130.990 55.955 ;
        RECT 130.240 55.495 130.990 55.665 ;
        RECT 131.630 55.665 131.885 55.955 ;
        RECT 132.055 55.835 132.385 56.215 ;
        RECT 131.630 55.495 132.380 55.665 ;
        RECT 130.240 54.505 130.470 55.495 ;
        RECT 130.640 54.675 130.990 55.325 ;
        RECT 131.630 54.675 131.980 55.325 ;
        RECT 132.150 54.505 132.380 55.495 ;
        RECT 130.240 54.335 130.990 54.505 ;
        RECT 130.235 53.665 130.565 54.165 ;
        RECT 130.735 53.835 130.990 54.335 ;
        RECT 131.630 54.335 132.380 54.505 ;
        RECT 131.630 53.835 131.885 54.335 ;
        RECT 132.055 53.665 132.385 54.165 ;
        RECT 132.555 53.835 132.725 55.955 ;
        RECT 133.085 55.855 133.415 56.215 ;
        RECT 133.585 55.825 134.080 55.995 ;
        RECT 134.285 55.825 135.140 55.995 ;
        RECT 132.955 54.635 133.415 55.685 ;
        RECT 132.895 53.850 133.220 54.635 ;
        RECT 133.585 54.465 133.755 55.825 ;
        RECT 133.925 54.915 134.275 55.535 ;
        RECT 134.445 55.315 134.800 55.535 ;
        RECT 134.445 54.725 134.615 55.315 ;
        RECT 134.970 55.115 135.140 55.825 ;
        RECT 136.015 55.755 136.345 56.215 ;
        RECT 136.555 55.855 136.905 56.025 ;
        RECT 135.345 55.285 136.135 55.535 ;
        RECT 136.555 55.465 136.815 55.855 ;
        RECT 137.125 55.765 138.075 56.045 ;
        RECT 138.245 55.775 138.435 56.215 ;
        RECT 138.605 55.835 139.675 56.005 ;
        RECT 136.305 55.115 136.475 55.295 ;
        RECT 133.585 54.295 133.980 54.465 ;
        RECT 134.150 54.335 134.615 54.725 ;
        RECT 134.785 54.945 136.475 55.115 ;
        RECT 133.810 54.165 133.980 54.295 ;
        RECT 134.785 54.165 134.955 54.945 ;
        RECT 136.645 54.775 136.815 55.465 ;
        RECT 135.315 54.605 136.815 54.775 ;
        RECT 137.005 54.805 137.215 55.595 ;
        RECT 137.385 54.975 137.735 55.595 ;
        RECT 137.905 54.985 138.075 55.765 ;
        RECT 138.605 55.605 138.775 55.835 ;
        RECT 138.245 55.435 138.775 55.605 ;
        RECT 138.245 55.155 138.465 55.435 ;
        RECT 138.945 55.265 139.185 55.665 ;
        RECT 137.905 54.815 138.310 54.985 ;
        RECT 138.645 54.895 139.185 55.265 ;
        RECT 139.355 55.480 139.675 55.835 ;
        RECT 139.920 55.755 140.225 56.215 ;
        RECT 140.395 55.505 140.650 56.035 ;
        RECT 139.355 55.305 139.680 55.480 ;
        RECT 139.355 55.005 140.270 55.305 ;
        RECT 139.530 54.975 140.270 55.005 ;
        RECT 137.005 54.645 137.680 54.805 ;
        RECT 138.140 54.725 138.310 54.815 ;
        RECT 137.005 54.635 137.970 54.645 ;
        RECT 136.645 54.465 136.815 54.605 ;
        RECT 133.390 53.665 133.640 54.125 ;
        RECT 133.810 53.835 134.060 54.165 ;
        RECT 134.275 53.835 134.955 54.165 ;
        RECT 135.125 54.265 136.200 54.435 ;
        RECT 136.645 54.295 137.205 54.465 ;
        RECT 137.510 54.345 137.970 54.635 ;
        RECT 138.140 54.555 139.360 54.725 ;
        RECT 135.125 53.925 135.295 54.265 ;
        RECT 135.530 53.665 135.860 54.095 ;
        RECT 136.030 53.925 136.200 54.265 ;
        RECT 136.495 53.665 136.865 54.125 ;
        RECT 137.035 53.835 137.205 54.295 ;
        RECT 138.140 54.175 138.310 54.555 ;
        RECT 139.530 54.385 139.700 54.975 ;
        RECT 140.440 54.855 140.650 55.505 ;
        RECT 140.885 55.395 141.095 56.215 ;
        RECT 141.265 55.415 141.595 56.045 ;
        RECT 137.440 53.835 138.310 54.175 ;
        RECT 138.900 54.215 139.700 54.385 ;
        RECT 138.480 53.665 138.730 54.125 ;
        RECT 138.900 53.925 139.070 54.215 ;
        RECT 139.250 53.665 139.580 54.045 ;
        RECT 139.920 53.665 140.225 54.805 ;
        RECT 140.395 53.975 140.650 54.855 ;
        RECT 141.265 54.815 141.515 55.415 ;
        RECT 141.765 55.395 141.995 56.215 ;
        RECT 142.665 55.490 142.955 56.215 ;
        RECT 143.125 55.445 145.715 56.215 ;
        RECT 141.685 54.975 142.015 55.225 ;
        RECT 143.125 54.925 144.335 55.445 ;
        RECT 146.385 55.395 146.615 56.215 ;
        RECT 146.785 55.415 147.115 56.045 ;
        RECT 140.885 53.665 141.095 54.805 ;
        RECT 141.265 53.835 141.595 54.815 ;
        RECT 141.765 53.665 141.995 54.805 ;
        RECT 142.665 53.665 142.955 54.830 ;
        RECT 144.505 54.755 145.715 55.275 ;
        RECT 146.365 54.975 146.695 55.225 ;
        RECT 146.865 54.815 147.115 55.415 ;
        RECT 147.285 55.395 147.495 56.215 ;
        RECT 147.725 55.445 150.315 56.215 ;
        RECT 150.945 55.465 152.155 56.215 ;
        RECT 147.725 54.925 148.935 55.445 ;
        RECT 143.125 53.665 145.715 54.755 ;
        RECT 146.385 53.665 146.615 54.805 ;
        RECT 146.785 53.835 147.115 54.815 ;
        RECT 147.285 53.665 147.495 54.805 ;
        RECT 149.105 54.755 150.315 55.275 ;
        RECT 147.725 53.665 150.315 54.755 ;
        RECT 150.945 54.755 151.465 55.295 ;
        RECT 151.635 54.925 152.155 55.465 ;
        RECT 150.945 53.665 152.155 54.755 ;
        RECT 6.025 51.390 6.380 53.590 ;
        RECT 91.060 53.495 152.240 53.665 ;
        RECT 91.145 52.405 92.355 53.495 ;
        RECT 92.530 52.825 92.785 53.325 ;
        RECT 92.955 52.995 93.285 53.495 ;
        RECT 92.530 52.655 93.280 52.825 ;
        RECT 6.020 50.910 6.380 51.390 ;
        RECT 91.145 51.695 91.665 52.235 ;
        RECT 91.835 51.865 92.355 52.405 ;
        RECT 92.530 51.835 92.880 52.485 ;
        RECT 91.145 50.945 92.355 51.695 ;
        RECT 93.050 51.665 93.280 52.655 ;
        RECT 92.530 51.495 93.280 51.665 ;
        RECT 92.530 51.205 92.785 51.495 ;
        RECT 92.955 50.945 93.285 51.325 ;
        RECT 93.455 51.205 93.625 53.325 ;
        RECT 93.795 52.525 94.120 53.310 ;
        RECT 94.290 53.035 94.540 53.495 ;
        RECT 94.710 52.995 94.960 53.325 ;
        RECT 95.175 52.995 95.855 53.325 ;
        RECT 94.710 52.865 94.880 52.995 ;
        RECT 94.485 52.695 94.880 52.865 ;
        RECT 93.855 51.475 94.315 52.525 ;
        RECT 94.485 51.335 94.655 52.695 ;
        RECT 95.050 52.435 95.515 52.825 ;
        RECT 94.825 51.625 95.175 52.245 ;
        RECT 95.345 51.845 95.515 52.435 ;
        RECT 95.685 52.215 95.855 52.995 ;
        RECT 96.025 52.895 96.195 53.235 ;
        RECT 96.430 53.065 96.760 53.495 ;
        RECT 96.930 52.895 97.100 53.235 ;
        RECT 97.395 53.035 97.765 53.495 ;
        RECT 96.025 52.725 97.100 52.895 ;
        RECT 97.935 52.865 98.105 53.325 ;
        RECT 98.340 52.985 99.210 53.325 ;
        RECT 99.380 53.035 99.630 53.495 ;
        RECT 97.545 52.695 98.105 52.865 ;
        RECT 97.545 52.555 97.715 52.695 ;
        RECT 96.215 52.385 97.715 52.555 ;
        RECT 98.410 52.525 98.870 52.815 ;
        RECT 95.685 52.045 97.375 52.215 ;
        RECT 95.345 51.625 95.700 51.845 ;
        RECT 95.870 51.335 96.040 52.045 ;
        RECT 96.245 51.625 97.035 51.875 ;
        RECT 97.205 51.865 97.375 52.045 ;
        RECT 97.545 51.695 97.715 52.385 ;
        RECT 93.985 50.945 94.315 51.305 ;
        RECT 94.485 51.165 94.980 51.335 ;
        RECT 95.185 51.165 96.040 51.335 ;
        RECT 96.915 50.945 97.245 51.405 ;
        RECT 97.455 51.305 97.715 51.695 ;
        RECT 97.905 52.515 98.870 52.525 ;
        RECT 99.040 52.605 99.210 52.985 ;
        RECT 99.800 52.945 99.970 53.235 ;
        RECT 100.150 53.115 100.480 53.495 ;
        RECT 99.800 52.775 100.600 52.945 ;
        RECT 97.905 52.355 98.580 52.515 ;
        RECT 99.040 52.435 100.260 52.605 ;
        RECT 97.905 51.565 98.115 52.355 ;
        RECT 99.040 52.345 99.210 52.435 ;
        RECT 98.285 51.565 98.635 52.185 ;
        RECT 98.805 52.175 99.210 52.345 ;
        RECT 98.805 51.395 98.975 52.175 ;
        RECT 99.145 51.725 99.365 52.005 ;
        RECT 99.545 51.895 100.085 52.265 ;
        RECT 100.430 52.185 100.600 52.775 ;
        RECT 100.820 52.355 101.125 53.495 ;
        RECT 101.295 52.305 101.550 53.185 ;
        RECT 101.785 52.355 101.995 53.495 ;
        RECT 100.430 52.155 101.170 52.185 ;
        RECT 99.145 51.555 99.675 51.725 ;
        RECT 97.455 51.135 97.805 51.305 ;
        RECT 98.025 51.115 98.975 51.395 ;
        RECT 99.145 50.945 99.335 51.385 ;
        RECT 99.505 51.325 99.675 51.555 ;
        RECT 99.845 51.495 100.085 51.895 ;
        RECT 100.255 51.855 101.170 52.155 ;
        RECT 100.255 51.680 100.580 51.855 ;
        RECT 100.255 51.325 100.575 51.680 ;
        RECT 101.340 51.655 101.550 52.305 ;
        RECT 102.165 52.345 102.495 53.325 ;
        RECT 102.665 52.355 102.895 53.495 ;
        RECT 99.505 51.155 100.575 51.325 ;
        RECT 100.820 50.945 101.125 51.405 ;
        RECT 101.295 51.125 101.550 51.655 ;
        RECT 101.785 50.945 101.995 51.765 ;
        RECT 102.165 51.745 102.415 52.345 ;
        RECT 104.025 52.330 104.315 53.495 ;
        RECT 104.485 52.405 106.155 53.495 ;
        RECT 102.585 51.935 102.915 52.185 ;
        RECT 102.165 51.115 102.495 51.745 ;
        RECT 102.665 50.945 102.895 51.765 ;
        RECT 104.485 51.715 105.235 52.235 ;
        RECT 105.405 51.885 106.155 52.405 ;
        RECT 106.510 52.525 106.900 52.700 ;
        RECT 107.385 52.695 107.715 53.495 ;
        RECT 107.885 52.705 108.420 53.325 ;
        RECT 106.510 52.355 107.935 52.525 ;
        RECT 104.025 50.945 104.315 51.670 ;
        RECT 104.485 50.945 106.155 51.715 ;
        RECT 106.385 51.625 106.740 52.185 ;
        RECT 106.910 51.455 107.080 52.355 ;
        RECT 107.250 51.625 107.515 52.185 ;
        RECT 107.765 51.855 107.935 52.355 ;
        RECT 108.105 51.685 108.420 52.705 ;
        RECT 106.490 50.945 106.730 51.455 ;
        RECT 106.910 51.125 107.190 51.455 ;
        RECT 107.420 50.945 107.635 51.455 ;
        RECT 107.805 51.115 108.420 51.685 ;
        RECT 109.085 52.420 109.355 53.325 ;
        RECT 109.525 52.735 109.855 53.495 ;
        RECT 110.035 52.565 110.205 53.325 ;
        RECT 109.085 51.620 109.255 52.420 ;
        RECT 109.540 52.395 110.205 52.565 ;
        RECT 111.110 52.525 111.500 52.700 ;
        RECT 111.985 52.695 112.315 53.495 ;
        RECT 112.485 52.705 113.020 53.325 ;
        RECT 109.540 52.250 109.710 52.395 ;
        RECT 111.110 52.355 112.535 52.525 ;
        RECT 109.425 51.920 109.710 52.250 ;
        RECT 109.540 51.665 109.710 51.920 ;
        RECT 109.945 51.845 110.275 52.215 ;
        RECT 109.085 51.115 109.345 51.620 ;
        RECT 109.540 51.495 110.205 51.665 ;
        RECT 110.985 51.625 111.340 52.185 ;
        RECT 109.525 50.945 109.855 51.325 ;
        RECT 110.035 51.115 110.205 51.495 ;
        RECT 111.510 51.455 111.680 52.355 ;
        RECT 111.850 51.625 112.115 52.185 ;
        RECT 112.365 51.855 112.535 52.355 ;
        RECT 112.705 51.685 113.020 52.705 ;
        RECT 113.230 52.825 113.485 53.325 ;
        RECT 113.655 52.995 113.985 53.495 ;
        RECT 113.230 52.655 113.980 52.825 ;
        RECT 113.230 51.835 113.580 52.485 ;
        RECT 111.090 50.945 111.330 51.455 ;
        RECT 111.510 51.125 111.790 51.455 ;
        RECT 112.020 50.945 112.235 51.455 ;
        RECT 112.405 51.115 113.020 51.685 ;
        RECT 113.750 51.665 113.980 52.655 ;
        RECT 113.230 51.495 113.980 51.665 ;
        RECT 113.230 51.205 113.485 51.495 ;
        RECT 113.655 50.945 113.985 51.325 ;
        RECT 114.155 51.205 114.325 53.325 ;
        RECT 114.495 52.525 114.820 53.310 ;
        RECT 114.990 53.035 115.240 53.495 ;
        RECT 115.410 52.995 115.660 53.325 ;
        RECT 115.875 52.995 116.555 53.325 ;
        RECT 115.410 52.865 115.580 52.995 ;
        RECT 115.185 52.695 115.580 52.865 ;
        RECT 114.555 51.475 115.015 52.525 ;
        RECT 115.185 51.335 115.355 52.695 ;
        RECT 115.750 52.435 116.215 52.825 ;
        RECT 115.525 51.625 115.875 52.245 ;
        RECT 116.045 51.845 116.215 52.435 ;
        RECT 116.385 52.215 116.555 52.995 ;
        RECT 116.725 52.895 116.895 53.235 ;
        RECT 117.130 53.065 117.460 53.495 ;
        RECT 117.630 52.895 117.800 53.235 ;
        RECT 118.095 53.035 118.465 53.495 ;
        RECT 116.725 52.725 117.800 52.895 ;
        RECT 118.635 52.865 118.805 53.325 ;
        RECT 119.040 52.985 119.910 53.325 ;
        RECT 120.080 53.035 120.330 53.495 ;
        RECT 118.245 52.695 118.805 52.865 ;
        RECT 118.245 52.555 118.415 52.695 ;
        RECT 116.915 52.385 118.415 52.555 ;
        RECT 119.110 52.525 119.570 52.815 ;
        RECT 116.385 52.045 118.075 52.215 ;
        RECT 116.045 51.625 116.400 51.845 ;
        RECT 116.570 51.335 116.740 52.045 ;
        RECT 116.945 51.625 117.735 51.875 ;
        RECT 117.905 51.865 118.075 52.045 ;
        RECT 118.245 51.695 118.415 52.385 ;
        RECT 114.685 50.945 115.015 51.305 ;
        RECT 115.185 51.165 115.680 51.335 ;
        RECT 115.885 51.165 116.740 51.335 ;
        RECT 117.615 50.945 117.945 51.405 ;
        RECT 118.155 51.305 118.415 51.695 ;
        RECT 118.605 52.515 119.570 52.525 ;
        RECT 119.740 52.605 119.910 52.985 ;
        RECT 120.500 52.945 120.670 53.235 ;
        RECT 120.850 53.115 121.180 53.495 ;
        RECT 120.500 52.775 121.300 52.945 ;
        RECT 118.605 52.355 119.280 52.515 ;
        RECT 119.740 52.435 120.960 52.605 ;
        RECT 118.605 51.565 118.815 52.355 ;
        RECT 119.740 52.345 119.910 52.435 ;
        RECT 118.985 51.565 119.335 52.185 ;
        RECT 119.505 52.175 119.910 52.345 ;
        RECT 119.505 51.395 119.675 52.175 ;
        RECT 119.845 51.725 120.065 52.005 ;
        RECT 120.245 51.895 120.785 52.265 ;
        RECT 121.130 52.185 121.300 52.775 ;
        RECT 121.520 52.355 121.825 53.495 ;
        RECT 121.995 52.305 122.250 53.185 ;
        RECT 123.545 52.825 123.825 53.495 ;
        RECT 123.995 52.605 124.295 53.155 ;
        RECT 124.495 52.775 124.825 53.495 ;
        RECT 125.015 52.775 125.475 53.325 ;
        RECT 125.645 52.985 125.905 53.495 ;
        RECT 121.130 52.155 121.870 52.185 ;
        RECT 119.845 51.555 120.375 51.725 ;
        RECT 118.155 51.135 118.505 51.305 ;
        RECT 118.725 51.115 119.675 51.395 ;
        RECT 119.845 50.945 120.035 51.385 ;
        RECT 120.205 51.325 120.375 51.555 ;
        RECT 120.545 51.495 120.785 51.895 ;
        RECT 120.955 51.855 121.870 52.155 ;
        RECT 120.955 51.680 121.280 51.855 ;
        RECT 120.955 51.325 121.275 51.680 ;
        RECT 122.040 51.655 122.250 52.305 ;
        RECT 123.360 52.185 123.625 52.545 ;
        RECT 123.995 52.435 124.935 52.605 ;
        RECT 124.765 52.185 124.935 52.435 ;
        RECT 123.360 51.935 124.035 52.185 ;
        RECT 124.255 51.935 124.595 52.185 ;
        RECT 124.765 51.855 125.055 52.185 ;
        RECT 124.765 51.765 124.935 51.855 ;
        RECT 120.205 51.155 121.275 51.325 ;
        RECT 121.520 50.945 121.825 51.405 ;
        RECT 121.995 51.125 122.250 51.655 ;
        RECT 123.545 51.575 124.935 51.765 ;
        RECT 123.545 51.215 123.875 51.575 ;
        RECT 125.225 51.405 125.475 52.775 ;
        RECT 125.645 51.935 125.985 52.815 ;
        RECT 126.155 52.105 126.325 53.325 ;
        RECT 126.565 52.990 127.180 53.495 ;
        RECT 126.565 52.455 126.815 52.820 ;
        RECT 126.985 52.815 127.180 52.990 ;
        RECT 127.350 52.985 127.825 53.325 ;
        RECT 127.995 52.950 128.210 53.495 ;
        RECT 126.985 52.625 127.315 52.815 ;
        RECT 127.535 52.455 128.250 52.750 ;
        RECT 128.420 52.625 128.695 53.325 ;
        RECT 126.565 52.285 128.355 52.455 ;
        RECT 126.155 51.855 126.950 52.105 ;
        RECT 126.155 51.765 126.405 51.855 ;
        RECT 124.495 50.945 124.745 51.405 ;
        RECT 124.915 51.115 125.475 51.405 ;
        RECT 125.645 50.945 125.905 51.765 ;
        RECT 126.075 51.345 126.405 51.765 ;
        RECT 127.120 51.430 127.375 52.285 ;
        RECT 126.585 51.165 127.375 51.430 ;
        RECT 127.545 51.585 127.955 52.105 ;
        RECT 128.125 51.855 128.355 52.285 ;
        RECT 128.525 51.595 128.695 52.625 ;
        RECT 129.785 52.330 130.075 53.495 ;
        RECT 131.165 52.625 131.440 53.325 ;
        RECT 131.650 52.950 131.865 53.495 ;
        RECT 132.035 52.985 132.510 53.325 ;
        RECT 132.680 52.990 133.295 53.495 ;
        RECT 132.680 52.815 132.875 52.990 ;
        RECT 127.545 51.165 127.745 51.585 ;
        RECT 127.935 50.945 128.265 51.405 ;
        RECT 128.435 51.115 128.695 51.595 ;
        RECT 129.785 50.945 130.075 51.670 ;
        RECT 131.165 51.595 131.335 52.625 ;
        RECT 131.610 52.455 132.325 52.750 ;
        RECT 132.545 52.625 132.875 52.815 ;
        RECT 133.045 52.455 133.295 52.820 ;
        RECT 131.505 52.285 133.295 52.455 ;
        RECT 131.505 51.855 131.735 52.285 ;
        RECT 131.165 51.115 131.425 51.595 ;
        RECT 131.905 51.585 132.315 52.105 ;
        RECT 131.595 50.945 131.925 51.405 ;
        RECT 132.115 51.165 132.315 51.585 ;
        RECT 132.485 51.430 132.740 52.285 ;
        RECT 133.535 52.105 133.705 53.325 ;
        RECT 133.955 52.985 134.215 53.495 ;
        RECT 132.910 51.855 133.705 52.105 ;
        RECT 133.875 51.935 134.215 52.815 ;
        RECT 134.385 52.625 134.660 53.325 ;
        RECT 134.830 52.950 135.085 53.495 ;
        RECT 135.255 52.985 135.735 53.325 ;
        RECT 135.910 52.940 136.515 53.495 ;
        RECT 136.685 52.985 136.945 53.495 ;
        RECT 135.900 52.840 136.515 52.940 ;
        RECT 135.900 52.815 136.085 52.840 ;
        RECT 133.455 51.765 133.705 51.855 ;
        RECT 132.485 51.165 133.275 51.430 ;
        RECT 133.455 51.345 133.785 51.765 ;
        RECT 133.955 50.945 134.215 51.765 ;
        RECT 134.385 51.595 134.555 52.625 ;
        RECT 134.830 52.495 135.585 52.745 ;
        RECT 135.755 52.570 136.085 52.815 ;
        RECT 134.830 52.460 135.600 52.495 ;
        RECT 134.830 52.450 135.615 52.460 ;
        RECT 134.725 52.435 135.620 52.450 ;
        RECT 134.725 52.420 135.640 52.435 ;
        RECT 134.725 52.410 135.660 52.420 ;
        RECT 134.725 52.400 135.685 52.410 ;
        RECT 134.725 52.370 135.755 52.400 ;
        RECT 134.725 52.340 135.775 52.370 ;
        RECT 134.725 52.310 135.795 52.340 ;
        RECT 134.725 52.285 135.825 52.310 ;
        RECT 134.725 52.250 135.860 52.285 ;
        RECT 134.725 52.245 135.890 52.250 ;
        RECT 134.725 51.850 134.955 52.245 ;
        RECT 135.500 52.240 135.890 52.245 ;
        RECT 135.525 52.230 135.890 52.240 ;
        RECT 135.540 52.225 135.890 52.230 ;
        RECT 135.555 52.220 135.890 52.225 ;
        RECT 136.255 52.220 136.515 52.670 ;
        RECT 135.555 52.215 136.515 52.220 ;
        RECT 135.565 52.205 136.515 52.215 ;
        RECT 135.575 52.200 136.515 52.205 ;
        RECT 135.585 52.190 136.515 52.200 ;
        RECT 135.590 52.180 136.515 52.190 ;
        RECT 135.595 52.175 136.515 52.180 ;
        RECT 135.605 52.160 136.515 52.175 ;
        RECT 135.610 52.145 136.515 52.160 ;
        RECT 135.620 52.120 136.515 52.145 ;
        RECT 135.125 51.650 135.455 52.075 ;
        RECT 134.385 51.115 134.645 51.595 ;
        RECT 134.815 50.945 135.065 51.485 ;
        RECT 135.235 51.165 135.455 51.650 ;
        RECT 135.625 52.050 136.515 52.120 ;
        RECT 135.625 51.325 135.795 52.050 ;
        RECT 136.685 51.935 137.025 52.815 ;
        RECT 137.195 52.105 137.365 53.325 ;
        RECT 137.605 52.990 138.220 53.495 ;
        RECT 137.605 52.455 137.855 52.820 ;
        RECT 138.025 52.815 138.220 52.990 ;
        RECT 138.390 52.985 138.865 53.325 ;
        RECT 139.035 52.950 139.250 53.495 ;
        RECT 138.025 52.625 138.355 52.815 ;
        RECT 138.575 52.455 139.290 52.750 ;
        RECT 139.460 52.625 139.735 53.325 ;
        RECT 137.605 52.285 139.395 52.455 ;
        RECT 135.965 51.495 136.515 51.880 ;
        RECT 137.195 51.855 137.990 52.105 ;
        RECT 137.195 51.765 137.445 51.855 ;
        RECT 135.625 51.155 136.515 51.325 ;
        RECT 136.685 50.945 136.945 51.765 ;
        RECT 137.115 51.345 137.445 51.765 ;
        RECT 138.160 51.430 138.415 52.285 ;
        RECT 137.625 51.165 138.415 51.430 ;
        RECT 138.585 51.585 138.995 52.105 ;
        RECT 139.165 51.855 139.395 52.285 ;
        RECT 139.565 51.595 139.735 52.625 ;
        RECT 139.995 52.565 140.165 53.325 ;
        RECT 140.345 52.735 140.675 53.495 ;
        RECT 139.995 52.395 140.660 52.565 ;
        RECT 140.845 52.420 141.115 53.325 ;
        RECT 141.290 52.825 141.545 53.325 ;
        RECT 141.715 52.995 142.045 53.495 ;
        RECT 141.290 52.655 142.040 52.825 ;
        RECT 140.490 52.250 140.660 52.395 ;
        RECT 139.925 51.845 140.255 52.215 ;
        RECT 140.490 51.920 140.775 52.250 ;
        RECT 140.490 51.665 140.660 51.920 ;
        RECT 138.585 51.165 138.785 51.585 ;
        RECT 138.975 50.945 139.305 51.405 ;
        RECT 139.475 51.115 139.735 51.595 ;
        RECT 139.995 51.495 140.660 51.665 ;
        RECT 140.945 51.620 141.115 52.420 ;
        RECT 141.290 51.835 141.640 52.485 ;
        RECT 141.810 51.665 142.040 52.655 ;
        RECT 139.995 51.115 140.165 51.495 ;
        RECT 140.345 50.945 140.675 51.325 ;
        RECT 140.855 51.115 141.115 51.620 ;
        RECT 141.290 51.495 142.040 51.665 ;
        RECT 141.290 51.205 141.545 51.495 ;
        RECT 141.715 50.945 142.045 51.325 ;
        RECT 142.215 51.205 142.385 53.325 ;
        RECT 142.555 52.525 142.880 53.310 ;
        RECT 143.050 53.035 143.300 53.495 ;
        RECT 143.470 52.995 143.720 53.325 ;
        RECT 143.935 52.995 144.615 53.325 ;
        RECT 143.470 52.865 143.640 52.995 ;
        RECT 143.245 52.695 143.640 52.865 ;
        RECT 142.615 51.475 143.075 52.525 ;
        RECT 143.245 51.335 143.415 52.695 ;
        RECT 143.810 52.435 144.275 52.825 ;
        RECT 143.585 51.625 143.935 52.245 ;
        RECT 144.105 51.845 144.275 52.435 ;
        RECT 144.445 52.215 144.615 52.995 ;
        RECT 144.785 52.895 144.955 53.235 ;
        RECT 145.190 53.065 145.520 53.495 ;
        RECT 145.690 52.895 145.860 53.235 ;
        RECT 146.155 53.035 146.525 53.495 ;
        RECT 144.785 52.725 145.860 52.895 ;
        RECT 146.695 52.865 146.865 53.325 ;
        RECT 147.100 52.985 147.970 53.325 ;
        RECT 148.140 53.035 148.390 53.495 ;
        RECT 146.305 52.695 146.865 52.865 ;
        RECT 146.305 52.555 146.475 52.695 ;
        RECT 144.975 52.385 146.475 52.555 ;
        RECT 147.170 52.525 147.630 52.815 ;
        RECT 144.445 52.045 146.135 52.215 ;
        RECT 144.105 51.625 144.460 51.845 ;
        RECT 144.630 51.335 144.800 52.045 ;
        RECT 145.005 51.625 145.795 51.875 ;
        RECT 145.965 51.865 146.135 52.045 ;
        RECT 146.305 51.695 146.475 52.385 ;
        RECT 142.745 50.945 143.075 51.305 ;
        RECT 143.245 51.165 143.740 51.335 ;
        RECT 143.945 51.165 144.800 51.335 ;
        RECT 145.675 50.945 146.005 51.405 ;
        RECT 146.215 51.305 146.475 51.695 ;
        RECT 146.665 52.515 147.630 52.525 ;
        RECT 147.800 52.605 147.970 52.985 ;
        RECT 148.560 52.945 148.730 53.235 ;
        RECT 148.910 53.115 149.240 53.495 ;
        RECT 148.560 52.775 149.360 52.945 ;
        RECT 146.665 52.355 147.340 52.515 ;
        RECT 147.800 52.435 149.020 52.605 ;
        RECT 146.665 51.565 146.875 52.355 ;
        RECT 147.800 52.345 147.970 52.435 ;
        RECT 147.045 51.565 147.395 52.185 ;
        RECT 147.565 52.175 147.970 52.345 ;
        RECT 147.565 51.395 147.735 52.175 ;
        RECT 147.905 51.725 148.125 52.005 ;
        RECT 148.305 51.895 148.845 52.265 ;
        RECT 149.190 52.185 149.360 52.775 ;
        RECT 149.580 52.355 149.885 53.495 ;
        RECT 150.055 52.305 150.310 53.185 ;
        RECT 149.190 52.155 149.930 52.185 ;
        RECT 147.905 51.555 148.435 51.725 ;
        RECT 146.215 51.135 146.565 51.305 ;
        RECT 146.785 51.115 147.735 51.395 ;
        RECT 147.905 50.945 148.095 51.385 ;
        RECT 148.265 51.325 148.435 51.555 ;
        RECT 148.605 51.495 148.845 51.895 ;
        RECT 149.015 51.855 149.930 52.155 ;
        RECT 149.015 51.680 149.340 51.855 ;
        RECT 149.015 51.325 149.335 51.680 ;
        RECT 150.100 51.655 150.310 52.305 ;
        RECT 150.945 52.405 152.155 53.495 ;
        RECT 150.945 51.865 151.465 52.405 ;
        RECT 151.635 51.695 152.155 52.235 ;
        RECT 148.265 51.155 149.335 51.325 ;
        RECT 149.580 50.945 149.885 51.405 ;
        RECT 150.055 51.125 150.310 51.655 ;
        RECT 150.945 50.945 152.155 51.695 ;
        RECT 6.025 46.455 6.380 50.910 ;
        RECT 91.060 50.775 152.240 50.945 ;
        RECT 91.145 50.025 92.355 50.775 ;
        RECT 91.145 49.485 91.665 50.025 ;
        RECT 92.525 50.005 96.035 50.775 ;
        RECT 96.205 50.025 97.415 50.775 ;
        RECT 97.585 50.100 97.845 50.605 ;
        RECT 98.025 50.395 98.355 50.775 ;
        RECT 98.535 50.225 98.705 50.605 ;
        RECT 91.835 49.315 92.355 49.855 ;
        RECT 92.525 49.485 94.175 50.005 ;
        RECT 94.345 49.315 96.035 49.835 ;
        RECT 96.205 49.485 96.725 50.025 ;
        RECT 96.895 49.315 97.415 49.855 ;
        RECT 91.145 48.225 92.355 49.315 ;
        RECT 92.525 48.225 96.035 49.315 ;
        RECT 96.205 48.225 97.415 49.315 ;
        RECT 97.585 49.300 97.755 50.100 ;
        RECT 98.040 50.055 98.705 50.225 ;
        RECT 98.040 49.800 98.210 50.055 ;
        RECT 99.025 49.955 99.235 50.775 ;
        RECT 99.405 49.975 99.735 50.605 ;
        RECT 97.925 49.470 98.210 49.800 ;
        RECT 98.445 49.505 98.775 49.875 ;
        RECT 98.040 49.325 98.210 49.470 ;
        RECT 99.405 49.375 99.655 49.975 ;
        RECT 99.905 49.955 100.135 50.775 ;
        RECT 100.345 50.005 102.015 50.775 ;
        RECT 102.385 50.145 102.715 50.505 ;
        RECT 103.335 50.315 103.585 50.775 ;
        RECT 103.755 50.315 104.315 50.605 ;
        RECT 99.825 49.535 100.155 49.785 ;
        RECT 100.345 49.485 101.095 50.005 ;
        RECT 102.385 49.955 103.775 50.145 ;
        RECT 103.605 49.865 103.775 49.955 ;
        RECT 97.585 48.395 97.855 49.300 ;
        RECT 98.040 49.155 98.705 49.325 ;
        RECT 98.025 48.225 98.355 48.985 ;
        RECT 98.535 48.395 98.705 49.155 ;
        RECT 99.025 48.225 99.235 49.365 ;
        RECT 99.405 48.395 99.735 49.375 ;
        RECT 99.905 48.225 100.135 49.365 ;
        RECT 101.265 49.315 102.015 49.835 ;
        RECT 100.345 48.225 102.015 49.315 ;
        RECT 102.200 49.535 102.875 49.785 ;
        RECT 103.095 49.535 103.435 49.785 ;
        RECT 103.605 49.535 103.895 49.865 ;
        RECT 102.200 49.175 102.465 49.535 ;
        RECT 103.605 49.285 103.775 49.535 ;
        RECT 102.835 49.115 103.775 49.285 ;
        RECT 102.385 48.225 102.665 48.895 ;
        RECT 102.835 48.565 103.135 49.115 ;
        RECT 104.065 48.945 104.315 50.315 ;
        RECT 103.335 48.225 103.665 48.945 ;
        RECT 103.855 48.395 104.315 48.945 ;
        RECT 104.945 50.125 105.205 50.605 ;
        RECT 105.375 50.235 105.625 50.775 ;
        RECT 104.945 49.095 105.115 50.125 ;
        RECT 105.795 50.070 106.015 50.555 ;
        RECT 105.285 49.475 105.515 49.870 ;
        RECT 105.685 49.645 106.015 50.070 ;
        RECT 106.185 50.395 107.075 50.565 ;
        RECT 106.185 49.670 106.355 50.395 ;
        RECT 107.250 50.225 107.505 50.515 ;
        RECT 107.675 50.395 108.005 50.775 ;
        RECT 106.525 49.840 107.075 50.225 ;
        RECT 107.250 50.055 108.000 50.225 ;
        RECT 106.185 49.600 107.075 49.670 ;
        RECT 106.180 49.575 107.075 49.600 ;
        RECT 106.170 49.560 107.075 49.575 ;
        RECT 106.165 49.545 107.075 49.560 ;
        RECT 106.155 49.540 107.075 49.545 ;
        RECT 106.150 49.530 107.075 49.540 ;
        RECT 106.145 49.520 107.075 49.530 ;
        RECT 106.135 49.515 107.075 49.520 ;
        RECT 106.125 49.505 107.075 49.515 ;
        RECT 106.115 49.500 107.075 49.505 ;
        RECT 106.115 49.495 106.450 49.500 ;
        RECT 106.100 49.490 106.450 49.495 ;
        RECT 106.085 49.480 106.450 49.490 ;
        RECT 106.060 49.475 106.450 49.480 ;
        RECT 105.285 49.470 106.450 49.475 ;
        RECT 105.285 49.435 106.420 49.470 ;
        RECT 105.285 49.410 106.385 49.435 ;
        RECT 105.285 49.380 106.355 49.410 ;
        RECT 105.285 49.350 106.335 49.380 ;
        RECT 105.285 49.320 106.315 49.350 ;
        RECT 105.285 49.310 106.245 49.320 ;
        RECT 105.285 49.300 106.220 49.310 ;
        RECT 105.285 49.285 106.200 49.300 ;
        RECT 105.285 49.270 106.180 49.285 ;
        RECT 105.390 49.260 106.175 49.270 ;
        RECT 105.390 49.225 106.160 49.260 ;
        RECT 104.945 48.395 105.220 49.095 ;
        RECT 105.390 48.975 106.145 49.225 ;
        RECT 106.315 48.905 106.645 49.150 ;
        RECT 106.815 49.050 107.075 49.500 ;
        RECT 107.250 49.235 107.600 49.885 ;
        RECT 107.770 49.065 108.000 50.055 ;
        RECT 106.460 48.880 106.645 48.905 ;
        RECT 107.250 48.895 108.000 49.065 ;
        RECT 106.460 48.780 107.075 48.880 ;
        RECT 105.390 48.225 105.645 48.770 ;
        RECT 105.815 48.395 106.295 48.735 ;
        RECT 106.470 48.225 107.075 48.780 ;
        RECT 107.250 48.395 107.505 48.895 ;
        RECT 107.675 48.225 108.005 48.725 ;
        RECT 108.175 48.395 108.345 50.515 ;
        RECT 108.705 50.415 109.035 50.775 ;
        RECT 109.205 50.385 109.700 50.555 ;
        RECT 109.905 50.385 110.760 50.555 ;
        RECT 108.575 49.195 109.035 50.245 ;
        RECT 108.515 48.410 108.840 49.195 ;
        RECT 109.205 49.025 109.375 50.385 ;
        RECT 109.545 49.475 109.895 50.095 ;
        RECT 110.065 49.875 110.420 50.095 ;
        RECT 110.065 49.285 110.235 49.875 ;
        RECT 110.590 49.675 110.760 50.385 ;
        RECT 111.635 50.315 111.965 50.775 ;
        RECT 112.175 50.415 112.525 50.585 ;
        RECT 110.965 49.845 111.755 50.095 ;
        RECT 112.175 50.025 112.435 50.415 ;
        RECT 112.745 50.325 113.695 50.605 ;
        RECT 113.865 50.335 114.055 50.775 ;
        RECT 114.225 50.395 115.295 50.565 ;
        RECT 111.925 49.675 112.095 49.855 ;
        RECT 109.205 48.855 109.600 49.025 ;
        RECT 109.770 48.895 110.235 49.285 ;
        RECT 110.405 49.505 112.095 49.675 ;
        RECT 109.430 48.725 109.600 48.855 ;
        RECT 110.405 48.725 110.575 49.505 ;
        RECT 112.265 49.335 112.435 50.025 ;
        RECT 110.935 49.165 112.435 49.335 ;
        RECT 112.625 49.365 112.835 50.155 ;
        RECT 113.005 49.535 113.355 50.155 ;
        RECT 113.525 49.545 113.695 50.325 ;
        RECT 114.225 50.165 114.395 50.395 ;
        RECT 113.865 49.995 114.395 50.165 ;
        RECT 113.865 49.715 114.085 49.995 ;
        RECT 114.565 49.825 114.805 50.225 ;
        RECT 113.525 49.375 113.930 49.545 ;
        RECT 114.265 49.455 114.805 49.825 ;
        RECT 114.975 50.040 115.295 50.395 ;
        RECT 115.540 50.315 115.845 50.775 ;
        RECT 116.015 50.065 116.265 50.595 ;
        RECT 114.975 49.865 115.300 50.040 ;
        RECT 114.975 49.565 115.890 49.865 ;
        RECT 115.150 49.535 115.890 49.565 ;
        RECT 112.625 49.205 113.300 49.365 ;
        RECT 113.760 49.285 113.930 49.375 ;
        RECT 112.625 49.195 113.590 49.205 ;
        RECT 112.265 49.025 112.435 49.165 ;
        RECT 109.010 48.225 109.260 48.685 ;
        RECT 109.430 48.395 109.680 48.725 ;
        RECT 109.895 48.395 110.575 48.725 ;
        RECT 110.745 48.825 111.820 48.995 ;
        RECT 112.265 48.855 112.825 49.025 ;
        RECT 113.130 48.905 113.590 49.195 ;
        RECT 113.760 49.115 114.980 49.285 ;
        RECT 110.745 48.485 110.915 48.825 ;
        RECT 111.150 48.225 111.480 48.655 ;
        RECT 111.650 48.485 111.820 48.825 ;
        RECT 112.115 48.225 112.485 48.685 ;
        RECT 112.655 48.395 112.825 48.855 ;
        RECT 113.760 48.735 113.930 49.115 ;
        RECT 115.150 48.945 115.320 49.535 ;
        RECT 116.060 49.415 116.265 50.065 ;
        RECT 116.435 50.020 116.685 50.775 ;
        RECT 116.905 50.050 117.195 50.775 ;
        RECT 117.365 50.230 122.710 50.775 ;
        RECT 113.060 48.395 113.930 48.735 ;
        RECT 114.520 48.775 115.320 48.945 ;
        RECT 114.100 48.225 114.350 48.685 ;
        RECT 114.520 48.485 114.690 48.775 ;
        RECT 114.870 48.225 115.200 48.605 ;
        RECT 115.540 48.225 115.845 49.365 ;
        RECT 116.015 48.535 116.265 49.415 ;
        RECT 118.950 49.400 119.290 50.230 ;
        RECT 122.885 50.005 126.395 50.775 ;
        RECT 126.730 50.265 126.970 50.775 ;
        RECT 127.150 50.265 127.430 50.595 ;
        RECT 127.660 50.265 127.875 50.775 ;
        RECT 116.435 48.225 116.685 49.365 ;
        RECT 116.905 48.225 117.195 49.390 ;
        RECT 120.770 48.660 121.120 49.910 ;
        RECT 122.885 49.485 124.535 50.005 ;
        RECT 124.705 49.315 126.395 49.835 ;
        RECT 126.625 49.535 126.980 50.095 ;
        RECT 127.150 49.365 127.320 50.265 ;
        RECT 127.490 49.535 127.755 50.095 ;
        RECT 128.045 50.035 128.660 50.605 ;
        RECT 128.005 49.365 128.175 49.865 ;
        RECT 117.365 48.225 122.710 48.660 ;
        RECT 122.885 48.225 126.395 49.315 ;
        RECT 126.750 49.195 128.175 49.365 ;
        RECT 126.750 49.020 127.140 49.195 ;
        RECT 127.625 48.225 127.955 49.025 ;
        RECT 128.345 49.015 128.660 50.035 ;
        RECT 128.865 50.005 131.455 50.775 ;
        RECT 132.170 50.275 132.665 50.605 ;
        RECT 128.865 49.485 130.075 50.005 ;
        RECT 130.245 49.315 131.455 49.835 ;
        RECT 128.125 48.395 128.660 49.015 ;
        RECT 128.865 48.225 131.455 49.315 ;
        RECT 132.085 48.785 132.325 50.095 ;
        RECT 132.495 49.365 132.665 50.275 ;
        RECT 132.885 49.535 133.235 50.500 ;
        RECT 133.415 49.535 133.715 50.505 ;
        RECT 133.895 49.535 134.175 50.505 ;
        RECT 134.355 49.975 134.625 50.775 ;
        RECT 134.795 50.055 135.135 50.565 ;
        RECT 135.470 50.265 135.710 50.775 ;
        RECT 135.890 50.265 136.170 50.595 ;
        RECT 136.400 50.265 136.615 50.775 ;
        RECT 134.370 49.535 134.700 49.785 ;
        RECT 134.370 49.365 134.685 49.535 ;
        RECT 132.495 49.195 134.685 49.365 ;
        RECT 132.090 48.225 132.425 48.605 ;
        RECT 132.595 48.395 132.845 49.195 ;
        RECT 133.065 48.225 133.395 48.945 ;
        RECT 133.580 48.395 133.830 49.195 ;
        RECT 134.295 48.225 134.625 49.025 ;
        RECT 134.875 48.655 135.135 50.055 ;
        RECT 135.365 49.535 135.720 50.095 ;
        RECT 135.890 49.365 136.060 50.265 ;
        RECT 136.230 49.535 136.495 50.095 ;
        RECT 136.785 50.035 137.400 50.605 ;
        RECT 136.745 49.365 136.915 49.865 ;
        RECT 135.490 49.195 136.915 49.365 ;
        RECT 135.490 49.020 135.880 49.195 ;
        RECT 134.795 48.395 135.135 48.655 ;
        RECT 136.365 48.225 136.695 49.025 ;
        RECT 137.085 49.015 137.400 50.035 ;
        RECT 137.605 50.005 141.115 50.775 ;
        RECT 141.285 50.025 142.495 50.775 ;
        RECT 142.665 50.050 142.955 50.775 ;
        RECT 137.605 49.485 139.255 50.005 ;
        RECT 139.425 49.315 141.115 49.835 ;
        RECT 141.285 49.485 141.805 50.025 ;
        RECT 143.125 50.005 145.715 50.775 ;
        RECT 146.345 50.035 146.605 50.605 ;
        RECT 146.775 50.375 147.160 50.775 ;
        RECT 147.330 50.205 147.585 50.605 ;
        RECT 146.775 50.035 147.585 50.205 ;
        RECT 147.775 50.035 148.020 50.605 ;
        RECT 148.190 50.375 148.575 50.775 ;
        RECT 148.745 50.205 149.000 50.605 ;
        RECT 148.190 50.035 149.000 50.205 ;
        RECT 149.190 50.035 149.615 50.605 ;
        RECT 149.785 50.375 150.170 50.775 ;
        RECT 150.340 50.205 150.775 50.605 ;
        RECT 149.785 50.035 150.775 50.205 ;
        RECT 141.975 49.315 142.495 49.855 ;
        RECT 143.125 49.485 144.335 50.005 ;
        RECT 136.865 48.395 137.400 49.015 ;
        RECT 137.605 48.225 141.115 49.315 ;
        RECT 141.285 48.225 142.495 49.315 ;
        RECT 142.665 48.225 142.955 49.390 ;
        RECT 144.505 49.315 145.715 49.835 ;
        RECT 143.125 48.225 145.715 49.315 ;
        RECT 146.345 49.365 146.530 50.035 ;
        RECT 146.775 49.865 147.125 50.035 ;
        RECT 147.775 49.865 147.945 50.035 ;
        RECT 148.190 49.865 148.540 50.035 ;
        RECT 149.190 49.865 149.540 50.035 ;
        RECT 149.785 49.865 150.120 50.035 ;
        RECT 150.945 50.025 152.155 50.775 ;
        RECT 146.700 49.535 147.125 49.865 ;
        RECT 146.345 48.395 146.605 49.365 ;
        RECT 146.775 49.015 147.125 49.535 ;
        RECT 147.295 49.365 147.945 49.865 ;
        RECT 148.115 49.535 148.540 49.865 ;
        RECT 147.295 49.185 148.020 49.365 ;
        RECT 146.775 48.820 147.585 49.015 ;
        RECT 146.775 48.225 147.160 48.650 ;
        RECT 147.330 48.395 147.585 48.820 ;
        RECT 147.775 48.395 148.020 49.185 ;
        RECT 148.190 49.015 148.540 49.535 ;
        RECT 148.710 49.365 149.540 49.865 ;
        RECT 149.710 49.535 150.120 49.865 ;
        RECT 148.710 49.185 149.615 49.365 ;
        RECT 148.190 48.820 149.020 49.015 ;
        RECT 148.190 48.225 148.575 48.650 ;
        RECT 148.745 48.395 149.020 48.820 ;
        RECT 149.190 48.395 149.615 49.185 ;
        RECT 149.785 48.990 150.120 49.535 ;
        RECT 150.290 49.160 150.775 49.865 ;
        RECT 150.945 49.315 151.465 49.855 ;
        RECT 151.635 49.485 152.155 50.025 ;
        RECT 149.785 48.820 150.775 48.990 ;
        RECT 149.785 48.225 150.170 48.650 ;
        RECT 150.340 48.395 150.775 48.820 ;
        RECT 150.945 48.225 152.155 49.315 ;
        RECT 91.060 48.055 152.240 48.225 ;
        RECT 91.145 46.965 92.355 48.055 ;
        RECT 92.990 47.385 93.245 47.885 ;
        RECT 93.415 47.555 93.745 48.055 ;
        RECT 92.990 47.215 93.740 47.385 ;
        RECT 6.030 44.420 6.380 46.455 ;
        RECT 91.145 46.255 91.665 46.795 ;
        RECT 91.835 46.425 92.355 46.965 ;
        RECT 92.990 46.395 93.340 47.045 ;
        RECT 91.145 45.505 92.355 46.255 ;
        RECT 93.510 46.225 93.740 47.215 ;
        RECT 92.990 46.055 93.740 46.225 ;
        RECT 92.990 45.765 93.245 46.055 ;
        RECT 93.415 45.505 93.745 45.885 ;
        RECT 93.915 45.765 94.085 47.885 ;
        RECT 94.255 47.085 94.580 47.870 ;
        RECT 94.750 47.595 95.000 48.055 ;
        RECT 95.170 47.555 95.420 47.885 ;
        RECT 95.635 47.555 96.315 47.885 ;
        RECT 95.170 47.425 95.340 47.555 ;
        RECT 94.945 47.255 95.340 47.425 ;
        RECT 94.315 46.035 94.775 47.085 ;
        RECT 94.945 45.895 95.115 47.255 ;
        RECT 95.510 46.995 95.975 47.385 ;
        RECT 95.285 46.185 95.635 46.805 ;
        RECT 95.805 46.405 95.975 46.995 ;
        RECT 96.145 46.775 96.315 47.555 ;
        RECT 96.485 47.455 96.655 47.795 ;
        RECT 96.890 47.625 97.220 48.055 ;
        RECT 97.390 47.455 97.560 47.795 ;
        RECT 97.855 47.595 98.225 48.055 ;
        RECT 96.485 47.285 97.560 47.455 ;
        RECT 98.395 47.425 98.565 47.885 ;
        RECT 98.800 47.545 99.670 47.885 ;
        RECT 99.840 47.595 100.090 48.055 ;
        RECT 98.005 47.255 98.565 47.425 ;
        RECT 98.005 47.115 98.175 47.255 ;
        RECT 96.675 46.945 98.175 47.115 ;
        RECT 98.870 47.085 99.330 47.375 ;
        RECT 96.145 46.605 97.835 46.775 ;
        RECT 95.805 46.185 96.160 46.405 ;
        RECT 96.330 45.895 96.500 46.605 ;
        RECT 96.705 46.185 97.495 46.435 ;
        RECT 97.665 46.425 97.835 46.605 ;
        RECT 98.005 46.255 98.175 46.945 ;
        RECT 94.445 45.505 94.775 45.865 ;
        RECT 94.945 45.725 95.440 45.895 ;
        RECT 95.645 45.725 96.500 45.895 ;
        RECT 97.375 45.505 97.705 45.965 ;
        RECT 97.915 45.865 98.175 46.255 ;
        RECT 98.365 47.075 99.330 47.085 ;
        RECT 99.500 47.165 99.670 47.545 ;
        RECT 100.260 47.505 100.430 47.795 ;
        RECT 100.610 47.675 100.940 48.055 ;
        RECT 100.260 47.335 101.060 47.505 ;
        RECT 98.365 46.915 99.040 47.075 ;
        RECT 99.500 46.995 100.720 47.165 ;
        RECT 98.365 46.125 98.575 46.915 ;
        RECT 99.500 46.905 99.670 46.995 ;
        RECT 98.745 46.125 99.095 46.745 ;
        RECT 99.265 46.735 99.670 46.905 ;
        RECT 99.265 45.955 99.435 46.735 ;
        RECT 99.605 46.285 99.825 46.565 ;
        RECT 100.005 46.455 100.545 46.825 ;
        RECT 100.890 46.745 101.060 47.335 ;
        RECT 101.280 46.915 101.585 48.055 ;
        RECT 101.755 46.865 102.005 47.745 ;
        RECT 102.175 46.915 102.425 48.055 ;
        RECT 102.645 46.965 103.855 48.055 ;
        RECT 100.890 46.715 101.630 46.745 ;
        RECT 99.605 46.115 100.135 46.285 ;
        RECT 97.915 45.695 98.265 45.865 ;
        RECT 98.485 45.675 99.435 45.955 ;
        RECT 99.605 45.505 99.795 45.945 ;
        RECT 99.965 45.885 100.135 46.115 ;
        RECT 100.305 46.055 100.545 46.455 ;
        RECT 100.715 46.415 101.630 46.715 ;
        RECT 100.715 46.240 101.040 46.415 ;
        RECT 100.715 45.885 101.035 46.240 ;
        RECT 101.800 46.215 102.005 46.865 ;
        RECT 99.965 45.715 101.035 45.885 ;
        RECT 101.280 45.505 101.585 45.965 ;
        RECT 101.755 45.685 102.005 46.215 ;
        RECT 102.175 45.505 102.425 46.260 ;
        RECT 102.645 46.255 103.165 46.795 ;
        RECT 103.335 46.425 103.855 46.965 ;
        RECT 104.025 46.890 104.315 48.055 ;
        RECT 105.405 47.545 105.665 48.055 ;
        RECT 105.405 46.495 105.745 47.375 ;
        RECT 105.915 46.665 106.085 47.885 ;
        RECT 106.325 47.550 106.940 48.055 ;
        RECT 106.325 47.015 106.575 47.380 ;
        RECT 106.745 47.375 106.940 47.550 ;
        RECT 107.110 47.545 107.585 47.885 ;
        RECT 107.755 47.510 107.970 48.055 ;
        RECT 106.745 47.185 107.075 47.375 ;
        RECT 107.295 47.015 108.010 47.310 ;
        RECT 108.180 47.185 108.455 47.885 ;
        RECT 108.715 47.310 108.985 48.055 ;
        RECT 109.615 48.050 115.890 48.055 ;
        RECT 106.325 46.845 108.115 47.015 ;
        RECT 105.915 46.415 106.710 46.665 ;
        RECT 105.915 46.325 106.165 46.415 ;
        RECT 102.645 45.505 103.855 46.255 ;
        RECT 104.025 45.505 104.315 46.230 ;
        RECT 105.405 45.505 105.665 46.325 ;
        RECT 105.835 45.905 106.165 46.325 ;
        RECT 106.880 45.990 107.135 46.845 ;
        RECT 106.345 45.725 107.135 45.990 ;
        RECT 107.305 46.145 107.715 46.665 ;
        RECT 107.885 46.415 108.115 46.845 ;
        RECT 108.285 46.155 108.455 47.185 ;
        RECT 109.155 47.140 109.445 47.880 ;
        RECT 109.615 47.325 109.870 48.050 ;
        RECT 110.055 47.155 110.315 47.880 ;
        RECT 110.485 47.325 110.730 48.050 ;
        RECT 110.915 47.155 111.175 47.880 ;
        RECT 111.345 47.325 111.590 48.050 ;
        RECT 111.775 47.155 112.035 47.880 ;
        RECT 112.205 47.325 112.450 48.050 ;
        RECT 112.620 47.155 112.880 47.880 ;
        RECT 113.050 47.325 113.310 48.050 ;
        RECT 113.480 47.155 113.740 47.880 ;
        RECT 113.910 47.325 114.170 48.050 ;
        RECT 114.340 47.155 114.600 47.880 ;
        RECT 114.770 47.325 115.030 48.050 ;
        RECT 115.200 47.155 115.460 47.880 ;
        RECT 115.630 47.255 115.890 48.050 ;
        RECT 110.055 47.140 115.460 47.155 ;
        RECT 108.715 46.915 115.460 47.140 ;
        RECT 108.715 46.325 109.880 46.915 ;
        RECT 116.060 46.745 116.310 47.880 ;
        RECT 116.490 47.245 116.750 48.055 ;
        RECT 116.925 46.745 117.170 47.885 ;
        RECT 117.350 47.245 117.645 48.055 ;
        RECT 117.830 46.865 118.085 47.745 ;
        RECT 118.255 46.915 118.560 48.055 ;
        RECT 118.900 47.675 119.230 48.055 ;
        RECT 119.410 47.505 119.580 47.795 ;
        RECT 119.750 47.595 120.000 48.055 ;
        RECT 118.780 47.335 119.580 47.505 ;
        RECT 120.170 47.545 121.040 47.885 ;
        RECT 110.050 46.495 117.170 46.745 ;
        RECT 108.715 46.155 115.460 46.325 ;
        RECT 107.305 45.725 107.505 46.145 ;
        RECT 107.695 45.505 108.025 45.965 ;
        RECT 108.195 45.675 108.455 46.155 ;
        RECT 108.715 45.505 109.015 45.985 ;
        RECT 109.185 45.700 109.445 46.155 ;
        RECT 109.615 45.505 109.875 45.985 ;
        RECT 110.055 45.700 110.315 46.155 ;
        RECT 110.485 45.505 110.735 45.985 ;
        RECT 110.915 45.700 111.175 46.155 ;
        RECT 111.345 45.505 111.595 45.985 ;
        RECT 111.775 45.700 112.035 46.155 ;
        RECT 112.205 45.505 112.450 45.985 ;
        RECT 112.620 45.700 112.895 46.155 ;
        RECT 113.065 45.505 113.310 45.985 ;
        RECT 113.480 45.700 113.740 46.155 ;
        RECT 113.910 45.505 114.170 45.985 ;
        RECT 114.340 45.700 114.600 46.155 ;
        RECT 114.770 45.505 115.030 45.985 ;
        RECT 115.200 45.700 115.460 46.155 ;
        RECT 115.630 45.505 115.890 46.065 ;
        RECT 116.060 45.685 116.310 46.495 ;
        RECT 116.490 45.505 116.750 46.030 ;
        RECT 116.920 45.685 117.170 46.495 ;
        RECT 117.340 46.185 117.655 46.745 ;
        RECT 117.830 46.215 118.040 46.865 ;
        RECT 118.780 46.745 118.950 47.335 ;
        RECT 120.170 47.165 120.340 47.545 ;
        RECT 121.275 47.425 121.445 47.885 ;
        RECT 121.615 47.595 121.985 48.055 ;
        RECT 122.280 47.455 122.450 47.795 ;
        RECT 122.620 47.625 122.950 48.055 ;
        RECT 123.185 47.455 123.355 47.795 ;
        RECT 119.120 46.995 120.340 47.165 ;
        RECT 120.510 47.085 120.970 47.375 ;
        RECT 121.275 47.255 121.835 47.425 ;
        RECT 122.280 47.285 123.355 47.455 ;
        RECT 123.525 47.555 124.205 47.885 ;
        RECT 124.420 47.555 124.670 47.885 ;
        RECT 124.840 47.595 125.090 48.055 ;
        RECT 121.665 47.115 121.835 47.255 ;
        RECT 120.510 47.075 121.475 47.085 ;
        RECT 120.170 46.905 120.340 46.995 ;
        RECT 120.800 46.915 121.475 47.075 ;
        RECT 118.210 46.715 118.950 46.745 ;
        RECT 118.210 46.415 119.125 46.715 ;
        RECT 118.800 46.240 119.125 46.415 ;
        RECT 117.350 45.505 117.655 46.015 ;
        RECT 117.830 45.685 118.085 46.215 ;
        RECT 118.255 45.505 118.560 45.965 ;
        RECT 118.805 45.885 119.125 46.240 ;
        RECT 119.295 46.455 119.835 46.825 ;
        RECT 120.170 46.735 120.575 46.905 ;
        RECT 119.295 46.055 119.535 46.455 ;
        RECT 120.015 46.285 120.235 46.565 ;
        RECT 119.705 46.115 120.235 46.285 ;
        RECT 119.705 45.885 119.875 46.115 ;
        RECT 120.405 45.955 120.575 46.735 ;
        RECT 120.745 46.125 121.095 46.745 ;
        RECT 121.265 46.125 121.475 46.915 ;
        RECT 121.665 46.945 123.165 47.115 ;
        RECT 121.665 46.255 121.835 46.945 ;
        RECT 123.525 46.775 123.695 47.555 ;
        RECT 124.500 47.425 124.670 47.555 ;
        RECT 122.005 46.605 123.695 46.775 ;
        RECT 123.865 46.995 124.330 47.385 ;
        RECT 124.500 47.255 124.895 47.425 ;
        RECT 122.005 46.425 122.175 46.605 ;
        RECT 118.805 45.715 119.875 45.885 ;
        RECT 120.045 45.505 120.235 45.945 ;
        RECT 120.405 45.675 121.355 45.955 ;
        RECT 121.665 45.865 121.925 46.255 ;
        RECT 122.345 46.185 123.135 46.435 ;
        RECT 121.575 45.695 121.925 45.865 ;
        RECT 122.135 45.505 122.465 45.965 ;
        RECT 123.340 45.895 123.510 46.605 ;
        RECT 123.865 46.405 124.035 46.995 ;
        RECT 123.680 46.185 124.035 46.405 ;
        RECT 124.205 46.185 124.555 46.805 ;
        RECT 124.725 45.895 124.895 47.255 ;
        RECT 125.260 47.085 125.585 47.870 ;
        RECT 125.065 46.035 125.525 47.085 ;
        RECT 123.340 45.725 124.195 45.895 ;
        RECT 124.400 45.725 124.895 45.895 ;
        RECT 125.065 45.505 125.395 45.865 ;
        RECT 125.755 45.765 125.925 47.885 ;
        RECT 126.095 47.555 126.425 48.055 ;
        RECT 126.595 47.385 126.850 47.885 ;
        RECT 126.100 47.215 126.850 47.385 ;
        RECT 126.100 46.225 126.330 47.215 ;
        RECT 126.500 46.395 126.850 47.045 ;
        RECT 127.065 46.915 127.295 48.055 ;
        RECT 127.465 46.905 127.795 47.885 ;
        RECT 127.965 46.915 128.175 48.055 ;
        RECT 128.405 46.965 129.615 48.055 ;
        RECT 127.045 46.495 127.375 46.745 ;
        RECT 126.100 46.055 126.850 46.225 ;
        RECT 126.095 45.505 126.425 45.885 ;
        RECT 126.595 45.765 126.850 46.055 ;
        RECT 127.065 45.505 127.295 46.325 ;
        RECT 127.545 46.305 127.795 46.905 ;
        RECT 127.465 45.675 127.795 46.305 ;
        RECT 127.965 45.505 128.175 46.325 ;
        RECT 128.405 46.255 128.925 46.795 ;
        RECT 129.095 46.425 129.615 46.965 ;
        RECT 129.785 46.890 130.075 48.055 ;
        RECT 130.245 47.620 135.590 48.055 ;
        RECT 135.765 47.620 141.110 48.055 ;
        RECT 141.285 47.620 146.630 48.055 ;
        RECT 128.405 45.505 129.615 46.255 ;
        RECT 129.785 45.505 130.075 46.230 ;
        RECT 131.830 46.050 132.170 46.880 ;
        RECT 133.650 46.370 134.000 47.620 ;
        RECT 137.350 46.050 137.690 46.880 ;
        RECT 139.170 46.370 139.520 47.620 ;
        RECT 142.870 46.050 143.210 46.880 ;
        RECT 144.690 46.370 145.040 47.620 ;
        RECT 146.805 46.965 150.315 48.055 ;
        RECT 146.805 46.275 148.455 46.795 ;
        RECT 148.625 46.445 150.315 46.965 ;
        RECT 150.945 46.965 152.155 48.055 ;
        RECT 150.945 46.425 151.465 46.965 ;
        RECT 130.245 45.505 135.590 46.050 ;
        RECT 135.765 45.505 141.110 46.050 ;
        RECT 141.285 45.505 146.630 46.050 ;
        RECT 146.805 45.505 150.315 46.275 ;
        RECT 151.635 46.255 152.155 46.795 ;
        RECT 150.945 45.505 152.155 46.255 ;
        RECT 91.060 45.335 152.240 45.505 ;
        RECT 91.145 44.585 92.355 45.335 ;
        RECT 91.145 44.045 91.665 44.585 ;
        RECT 92.525 44.565 96.035 45.335 ;
        RECT 96.295 44.685 96.465 45.165 ;
        RECT 96.645 44.855 96.885 45.335 ;
        RECT 97.135 44.685 97.305 45.165 ;
        RECT 97.475 44.855 97.805 45.335 ;
        RECT 97.975 44.685 98.145 45.165 ;
        RECT 91.835 43.875 92.355 44.415 ;
        RECT 92.525 44.045 94.175 44.565 ;
        RECT 96.295 44.515 96.930 44.685 ;
        RECT 97.135 44.515 98.145 44.685 ;
        RECT 98.315 44.535 98.645 45.335 ;
        RECT 99.425 44.685 99.685 45.165 ;
        RECT 99.855 44.875 100.185 45.335 ;
        RECT 100.375 44.695 100.575 45.115 ;
        RECT 94.345 43.875 96.035 44.395 ;
        RECT 96.760 44.345 96.930 44.515 ;
        RECT 97.645 44.485 98.145 44.515 ;
        RECT 96.210 44.105 96.590 44.345 ;
        RECT 96.760 44.175 97.260 44.345 ;
        RECT 96.760 43.935 96.930 44.175 ;
        RECT 97.650 43.975 98.145 44.485 ;
        RECT 6.030 41.370 6.380 43.420 ;
        RECT 91.145 42.785 92.355 43.875 ;
        RECT 92.525 42.785 96.035 43.875 ;
        RECT 96.215 43.765 96.930 43.935 ;
        RECT 97.135 43.805 98.145 43.975 ;
        RECT 96.215 42.955 96.545 43.765 ;
        RECT 96.715 42.785 96.955 43.585 ;
        RECT 97.135 42.955 97.305 43.805 ;
        RECT 97.475 42.785 97.805 43.585 ;
        RECT 97.975 42.955 98.145 43.805 ;
        RECT 98.315 42.785 98.645 43.935 ;
        RECT 99.425 43.655 99.595 44.685 ;
        RECT 99.765 43.995 99.995 44.425 ;
        RECT 100.165 44.175 100.575 44.695 ;
        RECT 100.745 44.850 101.535 45.115 ;
        RECT 100.745 43.995 101.000 44.850 ;
        RECT 101.715 44.515 102.045 44.935 ;
        RECT 102.215 44.515 102.475 45.335 ;
        RECT 102.645 44.565 104.315 45.335 ;
        RECT 104.520 44.595 105.135 45.165 ;
        RECT 105.305 44.825 105.520 45.335 ;
        RECT 105.750 44.825 106.030 45.155 ;
        RECT 106.210 44.825 106.450 45.335 ;
        RECT 101.715 44.425 101.965 44.515 ;
        RECT 101.170 44.175 101.965 44.425 ;
        RECT 99.765 43.825 101.555 43.995 ;
        RECT 99.425 42.955 99.700 43.655 ;
        RECT 99.870 43.530 100.585 43.825 ;
        RECT 100.805 43.465 101.135 43.655 ;
        RECT 99.910 42.785 100.125 43.330 ;
        RECT 100.295 42.955 100.770 43.295 ;
        RECT 100.940 43.290 101.135 43.465 ;
        RECT 101.305 43.460 101.555 43.825 ;
        RECT 100.940 42.785 101.555 43.290 ;
        RECT 101.795 42.955 101.965 44.175 ;
        RECT 102.135 43.465 102.475 44.345 ;
        RECT 102.645 44.045 103.395 44.565 ;
        RECT 103.565 43.875 104.315 44.395 ;
        RECT 102.215 42.785 102.475 43.295 ;
        RECT 102.645 42.785 104.315 43.875 ;
        RECT 104.520 43.575 104.835 44.595 ;
        RECT 105.005 43.925 105.175 44.425 ;
        RECT 105.425 44.095 105.690 44.655 ;
        RECT 105.860 43.925 106.030 44.825 ;
        RECT 106.200 44.095 106.555 44.655 ;
        RECT 106.785 44.565 110.295 45.335 ;
        RECT 110.465 44.615 110.805 45.125 ;
        RECT 106.785 44.045 108.435 44.565 ;
        RECT 105.005 43.755 106.430 43.925 ;
        RECT 108.605 43.875 110.295 44.395 ;
        RECT 104.520 42.955 105.055 43.575 ;
        RECT 105.225 42.785 105.555 43.585 ;
        RECT 106.040 43.580 106.430 43.755 ;
        RECT 106.785 42.785 110.295 43.875 ;
        RECT 110.465 43.215 110.725 44.615 ;
        RECT 110.975 44.535 111.245 45.335 ;
        RECT 110.900 44.095 111.230 44.345 ;
        RECT 111.425 44.095 111.705 45.065 ;
        RECT 111.885 44.095 112.185 45.065 ;
        RECT 112.365 44.095 112.715 45.060 ;
        RECT 112.935 44.835 113.430 45.165 ;
        RECT 110.915 43.925 111.230 44.095 ;
        RECT 112.935 43.925 113.105 44.835 ;
        RECT 110.915 43.755 113.105 43.925 ;
        RECT 110.465 42.955 110.805 43.215 ;
        RECT 110.975 42.785 111.305 43.585 ;
        RECT 111.770 42.955 112.020 43.755 ;
        RECT 112.205 42.785 112.535 43.505 ;
        RECT 112.755 42.955 113.005 43.755 ;
        RECT 113.275 43.345 113.515 44.655 ;
        RECT 113.745 44.515 113.955 45.335 ;
        RECT 114.125 44.535 114.455 45.165 ;
        RECT 114.125 43.935 114.375 44.535 ;
        RECT 114.625 44.515 114.855 45.335 ;
        RECT 115.065 44.565 116.735 45.335 ;
        RECT 116.905 44.610 117.195 45.335 ;
        RECT 117.365 44.565 120.875 45.335 ;
        RECT 121.045 44.585 122.255 45.335 ;
        RECT 122.540 44.705 122.825 45.165 ;
        RECT 122.995 44.875 123.265 45.335 ;
        RECT 114.545 44.095 114.875 44.345 ;
        RECT 115.065 44.045 115.815 44.565 ;
        RECT 113.175 42.785 113.510 43.165 ;
        RECT 113.745 42.785 113.955 43.925 ;
        RECT 114.125 42.955 114.455 43.935 ;
        RECT 114.625 42.785 114.855 43.925 ;
        RECT 115.985 43.875 116.735 44.395 ;
        RECT 117.365 44.045 119.015 44.565 ;
        RECT 115.065 42.785 116.735 43.875 ;
        RECT 116.905 42.785 117.195 43.950 ;
        RECT 119.185 43.875 120.875 44.395 ;
        RECT 121.045 44.045 121.565 44.585 ;
        RECT 122.540 44.535 123.495 44.705 ;
        RECT 121.735 43.875 122.255 44.415 ;
        RECT 117.365 42.785 120.875 43.875 ;
        RECT 121.045 42.785 122.255 43.875 ;
        RECT 122.425 43.805 123.115 44.365 ;
        RECT 123.285 43.635 123.495 44.535 ;
        RECT 122.540 43.415 123.495 43.635 ;
        RECT 123.665 44.365 124.065 45.165 ;
        RECT 124.255 44.705 124.535 45.165 ;
        RECT 125.055 44.875 125.380 45.335 ;
        RECT 124.255 44.535 125.380 44.705 ;
        RECT 125.550 44.595 125.935 45.165 ;
        RECT 126.115 44.615 126.445 45.335 ;
        RECT 126.990 44.935 128.605 45.105 ;
        RECT 128.775 44.935 129.105 45.335 ;
        RECT 128.435 44.765 128.605 44.935 ;
        RECT 129.275 44.860 129.610 45.120 ;
        RECT 124.930 44.425 125.380 44.535 ;
        RECT 123.665 43.805 124.760 44.365 ;
        RECT 124.930 44.095 125.485 44.425 ;
        RECT 122.540 42.955 122.825 43.415 ;
        RECT 122.995 42.785 123.265 43.245 ;
        RECT 123.665 42.955 124.065 43.805 ;
        RECT 124.930 43.635 125.380 44.095 ;
        RECT 125.655 43.925 125.935 44.595 ;
        RECT 126.170 44.095 126.520 44.425 ;
        RECT 126.830 44.095 127.250 44.760 ;
        RECT 127.420 44.315 127.710 44.755 ;
        RECT 127.900 44.315 128.170 44.755 ;
        RECT 128.435 44.595 128.995 44.765 ;
        RECT 128.825 44.425 128.995 44.595 ;
        RECT 128.380 44.315 128.630 44.425 ;
        RECT 127.420 44.145 127.715 44.315 ;
        RECT 127.900 44.145 128.175 44.315 ;
        RECT 128.380 44.145 128.635 44.315 ;
        RECT 127.420 44.095 127.710 44.145 ;
        RECT 127.900 44.095 128.170 44.145 ;
        RECT 128.380 44.095 128.630 44.145 ;
        RECT 128.825 44.095 129.130 44.425 ;
        RECT 126.170 43.975 126.375 44.095 ;
        RECT 124.255 43.415 125.380 43.635 ;
        RECT 124.255 42.955 124.535 43.415 ;
        RECT 125.055 42.785 125.380 43.245 ;
        RECT 125.550 42.955 125.935 43.925 ;
        RECT 126.165 43.805 126.375 43.975 ;
        RECT 128.825 43.925 128.995 44.095 ;
        RECT 126.625 43.755 128.995 43.925 ;
        RECT 126.195 43.125 126.365 43.625 ;
        RECT 126.625 43.295 126.795 43.755 ;
        RECT 127.025 43.375 128.450 43.545 ;
        RECT 127.025 43.125 127.355 43.375 ;
        RECT 126.195 42.955 127.355 43.125 ;
        RECT 127.580 42.785 127.910 43.205 ;
        RECT 128.165 42.955 128.450 43.375 ;
        RECT 128.695 42.785 129.025 43.585 ;
        RECT 129.355 43.505 129.610 44.860 ;
        RECT 129.785 44.585 130.995 45.335 ;
        RECT 129.785 44.045 130.305 44.585 ;
        RECT 131.225 44.515 131.435 45.335 ;
        RECT 131.605 44.535 131.935 45.165 ;
        RECT 130.475 43.875 130.995 44.415 ;
        RECT 131.605 43.935 131.855 44.535 ;
        RECT 132.105 44.515 132.335 45.335 ;
        RECT 133.525 44.515 133.735 45.335 ;
        RECT 133.905 44.535 134.235 45.165 ;
        RECT 132.025 44.095 132.355 44.345 ;
        RECT 133.905 43.935 134.155 44.535 ;
        RECT 134.405 44.515 134.635 45.335 ;
        RECT 134.845 44.565 136.515 45.335 ;
        RECT 134.325 44.095 134.655 44.345 ;
        RECT 134.845 44.045 135.595 44.565 ;
        RECT 136.685 44.535 136.995 45.335 ;
        RECT 137.200 44.535 137.895 45.165 ;
        RECT 138.230 44.825 138.470 45.335 ;
        RECT 138.650 44.825 138.930 45.155 ;
        RECT 139.160 44.825 139.375 45.335 ;
        RECT 129.275 42.995 129.610 43.505 ;
        RECT 129.785 42.785 130.995 43.875 ;
        RECT 131.225 42.785 131.435 43.925 ;
        RECT 131.605 42.955 131.935 43.935 ;
        RECT 132.105 42.785 132.335 43.925 ;
        RECT 133.525 42.785 133.735 43.925 ;
        RECT 133.905 42.955 134.235 43.935 ;
        RECT 134.405 42.785 134.635 43.925 ;
        RECT 135.765 43.875 136.515 44.395 ;
        RECT 136.695 44.095 137.030 44.365 ;
        RECT 137.200 43.935 137.370 44.535 ;
        RECT 137.540 44.095 137.875 44.345 ;
        RECT 138.125 44.095 138.480 44.655 ;
        RECT 134.845 42.785 136.515 43.875 ;
        RECT 136.685 42.785 136.965 43.925 ;
        RECT 137.135 42.955 137.465 43.935 ;
        RECT 138.650 43.925 138.820 44.825 ;
        RECT 138.990 44.095 139.255 44.655 ;
        RECT 139.545 44.595 140.160 45.165 ;
        RECT 140.365 44.955 141.255 45.125 ;
        RECT 139.505 43.925 139.675 44.425 ;
        RECT 137.635 42.785 137.895 43.925 ;
        RECT 138.250 43.755 139.675 43.925 ;
        RECT 138.250 43.580 138.640 43.755 ;
        RECT 139.125 42.785 139.455 43.585 ;
        RECT 139.845 43.575 140.160 44.595 ;
        RECT 140.365 44.400 140.915 44.785 ;
        RECT 141.085 44.230 141.255 44.955 ;
        RECT 140.365 44.160 141.255 44.230 ;
        RECT 141.425 44.630 141.645 45.115 ;
        RECT 141.815 44.795 142.065 45.335 ;
        RECT 142.235 44.685 142.495 45.165 ;
        RECT 141.425 44.205 141.755 44.630 ;
        RECT 140.365 44.135 141.260 44.160 ;
        RECT 140.365 44.120 141.270 44.135 ;
        RECT 140.365 44.105 141.275 44.120 ;
        RECT 140.365 44.100 141.285 44.105 ;
        RECT 140.365 44.090 141.290 44.100 ;
        RECT 140.365 44.080 141.295 44.090 ;
        RECT 140.365 44.075 141.305 44.080 ;
        RECT 140.365 44.065 141.315 44.075 ;
        RECT 140.365 44.060 141.325 44.065 ;
        RECT 140.365 43.610 140.625 44.060 ;
        RECT 140.990 44.055 141.325 44.060 ;
        RECT 140.990 44.050 141.340 44.055 ;
        RECT 140.990 44.040 141.355 44.050 ;
        RECT 140.990 44.035 141.380 44.040 ;
        RECT 141.925 44.035 142.155 44.430 ;
        RECT 140.990 44.030 142.155 44.035 ;
        RECT 141.020 43.995 142.155 44.030 ;
        RECT 141.055 43.970 142.155 43.995 ;
        RECT 141.085 43.940 142.155 43.970 ;
        RECT 141.105 43.910 142.155 43.940 ;
        RECT 141.125 43.880 142.155 43.910 ;
        RECT 141.195 43.870 142.155 43.880 ;
        RECT 141.220 43.860 142.155 43.870 ;
        RECT 141.240 43.845 142.155 43.860 ;
        RECT 141.260 43.830 142.155 43.845 ;
        RECT 141.265 43.820 142.050 43.830 ;
        RECT 141.280 43.785 142.050 43.820 ;
        RECT 139.625 42.955 140.160 43.575 ;
        RECT 140.795 43.465 141.125 43.710 ;
        RECT 141.295 43.535 142.050 43.785 ;
        RECT 142.325 43.655 142.495 44.685 ;
        RECT 142.665 44.610 142.955 45.335 ;
        RECT 143.125 44.660 143.385 45.165 ;
        RECT 143.565 44.955 143.895 45.335 ;
        RECT 144.075 44.785 144.245 45.165 ;
        RECT 140.795 43.440 140.980 43.465 ;
        RECT 140.365 43.340 140.980 43.440 ;
        RECT 140.365 42.785 140.970 43.340 ;
        RECT 141.145 42.955 141.625 43.295 ;
        RECT 141.795 42.785 142.050 43.330 ;
        RECT 142.220 42.955 142.495 43.655 ;
        RECT 142.665 42.785 142.955 43.950 ;
        RECT 143.125 43.860 143.295 44.660 ;
        RECT 143.580 44.615 144.245 44.785 ;
        RECT 143.580 44.360 143.750 44.615 ;
        RECT 144.505 44.565 146.175 45.335 ;
        RECT 143.465 44.030 143.750 44.360 ;
        RECT 143.985 44.065 144.315 44.435 ;
        RECT 144.505 44.045 145.255 44.565 ;
        RECT 146.385 44.515 146.615 45.335 ;
        RECT 146.785 44.535 147.115 45.165 ;
        RECT 143.580 43.885 143.750 44.030 ;
        RECT 143.125 42.955 143.395 43.860 ;
        RECT 143.580 43.715 144.245 43.885 ;
        RECT 145.425 43.875 146.175 44.395 ;
        RECT 146.365 44.095 146.695 44.345 ;
        RECT 146.865 43.935 147.115 44.535 ;
        RECT 147.285 44.515 147.495 45.335 ;
        RECT 147.725 44.565 150.315 45.335 ;
        RECT 150.945 44.585 152.155 45.335 ;
        RECT 147.725 44.045 148.935 44.565 ;
        RECT 143.565 42.785 143.895 43.545 ;
        RECT 144.075 42.955 144.245 43.715 ;
        RECT 144.505 42.785 146.175 43.875 ;
        RECT 146.385 42.785 146.615 43.925 ;
        RECT 146.785 42.955 147.115 43.935 ;
        RECT 147.285 42.785 147.495 43.925 ;
        RECT 149.105 43.875 150.315 44.395 ;
        RECT 147.725 42.785 150.315 43.875 ;
        RECT 150.945 43.875 151.465 44.415 ;
        RECT 151.635 44.045 152.155 44.585 ;
        RECT 150.945 42.785 152.155 43.875 ;
        RECT 91.060 42.615 152.240 42.785 ;
        RECT 91.145 41.525 92.355 42.615 ;
        RECT 6.025 41.260 6.380 41.370 ;
        RECT 6.025 34.100 6.375 41.260 ;
        RECT 91.145 40.815 91.665 41.355 ;
        RECT 91.835 40.985 92.355 41.525 ;
        RECT 92.615 41.685 92.785 42.445 ;
        RECT 92.965 41.855 93.295 42.615 ;
        RECT 92.615 41.515 93.280 41.685 ;
        RECT 93.465 41.540 93.735 42.445 ;
        RECT 93.110 41.370 93.280 41.515 ;
        RECT 92.545 40.965 92.875 41.335 ;
        RECT 93.110 41.040 93.395 41.370 ;
        RECT 91.145 40.065 92.355 40.815 ;
        RECT 93.110 40.785 93.280 41.040 ;
        RECT 92.615 40.615 93.280 40.785 ;
        RECT 93.565 40.740 93.735 41.540 ;
        RECT 93.905 41.525 97.415 42.615 ;
        RECT 97.585 41.525 98.795 42.615 ;
        RECT 92.615 40.235 92.785 40.615 ;
        RECT 92.965 40.065 93.295 40.445 ;
        RECT 93.475 40.235 93.735 40.740 ;
        RECT 93.905 40.835 95.555 41.355 ;
        RECT 95.725 41.005 97.415 41.525 ;
        RECT 93.905 40.065 97.415 40.835 ;
        RECT 97.585 40.815 98.105 41.355 ;
        RECT 98.275 40.985 98.795 41.525 ;
        RECT 98.975 41.635 99.305 42.445 ;
        RECT 99.475 41.815 99.715 42.615 ;
        RECT 98.975 41.465 99.690 41.635 ;
        RECT 98.970 41.055 99.350 41.295 ;
        RECT 99.520 41.225 99.690 41.465 ;
        RECT 99.895 41.595 100.065 42.445 ;
        RECT 100.235 41.815 100.565 42.615 ;
        RECT 100.735 41.595 100.905 42.445 ;
        RECT 99.895 41.425 100.905 41.595 ;
        RECT 101.075 41.465 101.405 42.615 ;
        RECT 101.725 41.525 103.395 42.615 ;
        RECT 99.520 41.055 100.020 41.225 ;
        RECT 99.520 40.885 99.690 41.055 ;
        RECT 100.410 40.885 100.905 41.425 ;
        RECT 97.585 40.065 98.795 40.815 ;
        RECT 99.055 40.715 99.690 40.885 ;
        RECT 99.895 40.715 100.905 40.885 ;
        RECT 99.055 40.235 99.225 40.715 ;
        RECT 99.405 40.065 99.645 40.545 ;
        RECT 99.895 40.235 100.065 40.715 ;
        RECT 100.235 40.065 100.565 40.545 ;
        RECT 100.735 40.235 100.905 40.715 ;
        RECT 101.075 40.065 101.405 40.865 ;
        RECT 101.725 40.835 102.475 41.355 ;
        RECT 102.645 41.005 103.395 41.525 ;
        RECT 104.025 41.450 104.315 42.615 ;
        RECT 104.485 42.180 109.830 42.615 ;
        RECT 110.005 42.180 115.350 42.615 ;
        RECT 115.525 42.180 120.870 42.615 ;
        RECT 121.045 42.180 126.390 42.615 ;
        RECT 101.725 40.065 103.395 40.835 ;
        RECT 104.025 40.065 104.315 40.790 ;
        RECT 106.070 40.610 106.410 41.440 ;
        RECT 107.890 40.930 108.240 42.180 ;
        RECT 111.590 40.610 111.930 41.440 ;
        RECT 113.410 40.930 113.760 42.180 ;
        RECT 117.110 40.610 117.450 41.440 ;
        RECT 118.930 40.930 119.280 42.180 ;
        RECT 122.630 40.610 122.970 41.440 ;
        RECT 124.450 40.930 124.800 42.180 ;
        RECT 126.565 41.525 129.155 42.615 ;
        RECT 126.565 40.835 127.775 41.355 ;
        RECT 127.945 41.005 129.155 41.525 ;
        RECT 129.785 41.450 130.075 42.615 ;
        RECT 130.245 42.180 135.590 42.615 ;
        RECT 104.485 40.065 109.830 40.610 ;
        RECT 110.005 40.065 115.350 40.610 ;
        RECT 115.525 40.065 120.870 40.610 ;
        RECT 121.045 40.065 126.390 40.610 ;
        RECT 126.565 40.065 129.155 40.835 ;
        RECT 129.785 40.065 130.075 40.790 ;
        RECT 131.830 40.610 132.170 41.440 ;
        RECT 133.650 40.930 134.000 42.180 ;
        RECT 135.765 41.525 138.355 42.615 ;
        RECT 135.765 40.835 136.975 41.355 ;
        RECT 137.145 41.005 138.355 41.525 ;
        RECT 138.995 41.645 139.325 42.430 ;
        RECT 138.995 41.475 139.675 41.645 ;
        RECT 139.855 41.475 140.185 42.615 ;
        RECT 141.290 41.945 141.545 42.445 ;
        RECT 141.715 42.115 142.045 42.615 ;
        RECT 141.290 41.775 142.040 41.945 ;
        RECT 138.985 41.055 139.335 41.305 ;
        RECT 139.505 40.875 139.675 41.475 ;
        RECT 139.845 41.055 140.195 41.305 ;
        RECT 141.290 40.955 141.640 41.605 ;
        RECT 130.245 40.065 135.590 40.610 ;
        RECT 135.765 40.065 138.355 40.835 ;
        RECT 139.005 40.065 139.245 40.875 ;
        RECT 139.415 40.235 139.745 40.875 ;
        RECT 139.915 40.065 140.185 40.875 ;
        RECT 141.810 40.785 142.040 41.775 ;
        RECT 141.290 40.615 142.040 40.785 ;
        RECT 141.290 40.325 141.545 40.615 ;
        RECT 141.715 40.065 142.045 40.445 ;
        RECT 142.215 40.325 142.385 42.445 ;
        RECT 142.555 41.645 142.880 42.430 ;
        RECT 143.050 42.155 143.300 42.615 ;
        RECT 143.470 42.115 143.720 42.445 ;
        RECT 143.935 42.115 144.615 42.445 ;
        RECT 143.470 41.985 143.640 42.115 ;
        RECT 143.245 41.815 143.640 41.985 ;
        RECT 142.615 40.595 143.075 41.645 ;
        RECT 143.245 40.455 143.415 41.815 ;
        RECT 143.810 41.555 144.275 41.945 ;
        RECT 143.585 40.745 143.935 41.365 ;
        RECT 144.105 40.965 144.275 41.555 ;
        RECT 144.445 41.335 144.615 42.115 ;
        RECT 144.785 42.015 144.955 42.355 ;
        RECT 145.190 42.185 145.520 42.615 ;
        RECT 145.690 42.015 145.860 42.355 ;
        RECT 146.155 42.155 146.525 42.615 ;
        RECT 144.785 41.845 145.860 42.015 ;
        RECT 146.695 41.985 146.865 42.445 ;
        RECT 147.100 42.105 147.970 42.445 ;
        RECT 148.140 42.155 148.390 42.615 ;
        RECT 146.305 41.815 146.865 41.985 ;
        RECT 146.305 41.675 146.475 41.815 ;
        RECT 144.975 41.505 146.475 41.675 ;
        RECT 147.170 41.645 147.630 41.935 ;
        RECT 144.445 41.165 146.135 41.335 ;
        RECT 144.105 40.745 144.460 40.965 ;
        RECT 144.630 40.455 144.800 41.165 ;
        RECT 145.005 40.745 145.795 40.995 ;
        RECT 145.965 40.985 146.135 41.165 ;
        RECT 146.305 40.815 146.475 41.505 ;
        RECT 142.745 40.065 143.075 40.425 ;
        RECT 143.245 40.285 143.740 40.455 ;
        RECT 143.945 40.285 144.800 40.455 ;
        RECT 145.675 40.065 146.005 40.525 ;
        RECT 146.215 40.425 146.475 40.815 ;
        RECT 146.665 41.635 147.630 41.645 ;
        RECT 147.800 41.725 147.970 42.105 ;
        RECT 148.560 42.065 148.730 42.355 ;
        RECT 148.910 42.235 149.240 42.615 ;
        RECT 148.560 41.895 149.360 42.065 ;
        RECT 146.665 41.475 147.340 41.635 ;
        RECT 147.800 41.555 149.020 41.725 ;
        RECT 146.665 40.685 146.875 41.475 ;
        RECT 147.800 41.465 147.970 41.555 ;
        RECT 147.045 40.685 147.395 41.305 ;
        RECT 147.565 41.295 147.970 41.465 ;
        RECT 147.565 40.515 147.735 41.295 ;
        RECT 147.905 40.845 148.125 41.125 ;
        RECT 148.305 41.015 148.845 41.385 ;
        RECT 149.190 41.305 149.360 41.895 ;
        RECT 149.580 41.475 149.885 42.615 ;
        RECT 150.055 41.425 150.310 42.305 ;
        RECT 149.190 41.275 149.930 41.305 ;
        RECT 147.905 40.675 148.435 40.845 ;
        RECT 146.215 40.255 146.565 40.425 ;
        RECT 146.785 40.235 147.735 40.515 ;
        RECT 147.905 40.065 148.095 40.505 ;
        RECT 148.265 40.445 148.435 40.675 ;
        RECT 148.605 40.615 148.845 41.015 ;
        RECT 149.015 40.975 149.930 41.275 ;
        RECT 149.015 40.800 149.340 40.975 ;
        RECT 149.015 40.445 149.335 40.800 ;
        RECT 150.100 40.775 150.310 41.425 ;
        RECT 150.945 41.525 152.155 42.615 ;
        RECT 150.945 40.985 151.465 41.525 ;
        RECT 151.635 40.815 152.155 41.355 ;
        RECT 148.265 40.275 149.335 40.445 ;
        RECT 149.580 40.065 149.885 40.525 ;
        RECT 150.055 40.245 150.310 40.775 ;
        RECT 150.945 40.065 152.155 40.815 ;
        RECT 91.060 39.895 152.240 40.065 ;
        RECT 91.145 39.145 92.355 39.895 ;
        RECT 91.145 38.605 91.665 39.145 ;
        RECT 92.525 39.125 96.035 39.895 ;
        RECT 96.670 39.390 97.005 39.895 ;
        RECT 97.175 39.325 97.415 39.700 ;
        RECT 97.695 39.565 97.865 39.710 ;
        RECT 97.695 39.370 98.070 39.565 ;
        RECT 98.430 39.400 98.825 39.895 ;
        RECT 91.835 38.435 92.355 38.975 ;
        RECT 92.525 38.605 94.175 39.125 ;
        RECT 94.345 38.435 96.035 38.955 ;
        RECT 91.145 37.345 92.355 38.435 ;
        RECT 92.525 37.345 96.035 38.435 ;
        RECT 96.725 38.365 97.025 39.215 ;
        RECT 97.195 39.175 97.415 39.325 ;
        RECT 97.195 38.845 97.730 39.175 ;
        RECT 97.900 39.035 98.070 39.370 ;
        RECT 98.995 39.205 99.235 39.725 ;
        RECT 97.195 38.195 97.430 38.845 ;
        RECT 97.900 38.675 98.885 39.035 ;
        RECT 96.755 37.965 97.430 38.195 ;
        RECT 97.600 38.655 98.885 38.675 ;
        RECT 97.600 38.505 98.460 38.655 ;
        RECT 96.755 37.535 96.925 37.965 ;
        RECT 97.095 37.345 97.425 37.795 ;
        RECT 97.600 37.560 97.885 38.505 ;
        RECT 99.060 38.400 99.235 39.205 ;
        RECT 99.910 39.245 100.220 39.715 ;
        RECT 100.390 39.415 101.125 39.895 ;
        RECT 101.295 39.325 101.465 39.675 ;
        RECT 101.635 39.495 102.015 39.895 ;
        RECT 99.910 39.075 100.645 39.245 ;
        RECT 101.295 39.155 102.035 39.325 ;
        RECT 102.205 39.220 102.475 39.565 ;
        RECT 100.395 38.985 100.645 39.075 ;
        RECT 101.865 38.985 102.035 39.155 ;
        RECT 99.890 38.655 100.225 38.905 ;
        RECT 100.395 38.655 101.135 38.985 ;
        RECT 101.865 38.655 102.095 38.985 ;
        RECT 98.060 38.025 98.755 38.335 ;
        RECT 98.065 37.345 98.750 37.815 ;
        RECT 98.930 37.615 99.235 38.400 ;
        RECT 99.890 37.345 100.145 38.485 ;
        RECT 100.395 38.095 100.565 38.655 ;
        RECT 101.865 38.485 102.035 38.655 ;
        RECT 102.305 38.485 102.475 39.220 ;
        RECT 102.645 39.145 103.855 39.895 ;
        RECT 104.030 39.390 104.365 39.895 ;
        RECT 104.535 39.325 104.775 39.700 ;
        RECT 105.055 39.565 105.225 39.710 ;
        RECT 105.055 39.370 105.430 39.565 ;
        RECT 105.790 39.400 106.185 39.895 ;
        RECT 102.645 38.605 103.165 39.145 ;
        RECT 100.790 38.315 102.035 38.485 ;
        RECT 100.790 38.065 101.210 38.315 ;
        RECT 100.340 37.565 101.535 37.895 ;
        RECT 101.715 37.345 101.995 38.145 ;
        RECT 102.205 37.515 102.475 38.485 ;
        RECT 103.335 38.435 103.855 38.975 ;
        RECT 102.645 37.345 103.855 38.435 ;
        RECT 104.085 38.365 104.385 39.215 ;
        RECT 104.555 39.175 104.775 39.325 ;
        RECT 104.555 38.845 105.090 39.175 ;
        RECT 105.260 39.035 105.430 39.370 ;
        RECT 106.355 39.205 106.595 39.725 ;
        RECT 104.555 38.195 104.790 38.845 ;
        RECT 105.260 38.675 106.245 39.035 ;
        RECT 104.115 37.965 104.790 38.195 ;
        RECT 104.960 38.655 106.245 38.675 ;
        RECT 104.960 38.505 105.820 38.655 ;
        RECT 104.115 37.535 104.285 37.965 ;
        RECT 104.455 37.345 104.785 37.795 ;
        RECT 104.960 37.560 105.245 38.505 ;
        RECT 106.420 38.400 106.595 39.205 ;
        RECT 106.785 39.145 107.995 39.895 ;
        RECT 108.165 39.285 108.505 39.700 ;
        RECT 108.675 39.455 108.845 39.895 ;
        RECT 109.015 39.505 110.265 39.685 ;
        RECT 109.015 39.285 109.345 39.505 ;
        RECT 110.535 39.435 110.705 39.895 ;
        RECT 106.785 38.605 107.305 39.145 ;
        RECT 108.165 39.115 109.345 39.285 ;
        RECT 109.515 39.265 109.880 39.335 ;
        RECT 109.515 39.085 110.765 39.265 ;
        RECT 107.475 38.435 107.995 38.975 ;
        RECT 108.165 38.705 108.630 38.905 ;
        RECT 108.805 38.655 109.135 38.905 ;
        RECT 109.305 38.875 109.770 38.905 ;
        RECT 109.305 38.705 109.775 38.875 ;
        RECT 109.305 38.655 109.770 38.705 ;
        RECT 109.965 38.655 110.320 38.905 ;
        RECT 108.805 38.535 108.985 38.655 ;
        RECT 105.420 38.025 106.115 38.335 ;
        RECT 105.425 37.345 106.110 37.815 ;
        RECT 106.290 37.615 106.595 38.400 ;
        RECT 106.785 37.345 107.995 38.435 ;
        RECT 108.165 37.345 108.485 38.525 ;
        RECT 108.655 38.365 108.985 38.535 ;
        RECT 110.490 38.485 110.765 39.085 ;
        RECT 108.655 37.575 108.855 38.365 ;
        RECT 109.155 38.275 110.765 38.485 ;
        RECT 109.155 38.175 109.565 38.275 ;
        RECT 109.180 37.515 109.565 38.175 ;
        RECT 109.960 37.345 110.745 38.105 ;
        RECT 110.935 37.515 111.215 39.615 ;
        RECT 111.405 39.205 111.645 39.725 ;
        RECT 111.815 39.400 112.210 39.895 ;
        RECT 112.775 39.565 112.945 39.710 ;
        RECT 112.570 39.370 112.945 39.565 ;
        RECT 111.405 38.400 111.580 39.205 ;
        RECT 112.570 39.035 112.740 39.370 ;
        RECT 113.225 39.325 113.465 39.700 ;
        RECT 113.635 39.390 113.970 39.895 ;
        RECT 114.150 39.365 114.440 39.715 ;
        RECT 114.635 39.535 114.965 39.895 ;
        RECT 115.135 39.365 115.365 39.670 ;
        RECT 113.225 39.175 113.445 39.325 ;
        RECT 111.755 38.675 112.740 39.035 ;
        RECT 112.910 38.845 113.445 39.175 ;
        RECT 111.755 38.655 113.040 38.675 ;
        RECT 112.180 38.505 113.040 38.655 ;
        RECT 111.405 37.615 111.710 38.400 ;
        RECT 111.885 38.025 112.580 38.335 ;
        RECT 111.890 37.345 112.575 37.815 ;
        RECT 112.755 37.560 113.040 38.505 ;
        RECT 113.210 38.195 113.445 38.845 ;
        RECT 113.615 38.365 113.915 39.215 ;
        RECT 114.150 39.195 115.365 39.365 ;
        RECT 115.555 39.025 115.725 39.590 ;
        RECT 116.905 39.170 117.195 39.895 ;
        RECT 114.210 38.875 114.470 38.985 ;
        RECT 114.205 38.705 114.470 38.875 ;
        RECT 114.210 38.655 114.470 38.705 ;
        RECT 114.650 38.655 115.035 38.985 ;
        RECT 115.205 38.855 115.725 39.025 ;
        RECT 117.365 39.125 119.035 39.895 ;
        RECT 119.205 39.155 119.645 39.715 ;
        RECT 119.815 39.155 120.265 39.895 ;
        RECT 120.435 39.325 120.605 39.725 ;
        RECT 120.775 39.495 121.195 39.895 ;
        RECT 121.365 39.325 121.595 39.725 ;
        RECT 120.435 39.155 121.595 39.325 ;
        RECT 121.765 39.155 122.255 39.725 ;
        RECT 113.210 37.965 113.885 38.195 ;
        RECT 113.215 37.345 113.545 37.795 ;
        RECT 113.715 37.535 113.885 37.965 ;
        RECT 114.150 37.345 114.470 38.485 ;
        RECT 114.650 37.605 114.845 38.655 ;
        RECT 115.205 38.475 115.375 38.855 ;
        RECT 115.025 38.195 115.375 38.475 ;
        RECT 115.565 38.325 115.810 38.685 ;
        RECT 117.365 38.605 118.115 39.125 ;
        RECT 115.025 37.515 115.355 38.195 ;
        RECT 115.555 37.345 115.810 38.145 ;
        RECT 116.905 37.345 117.195 38.510 ;
        RECT 118.285 38.435 119.035 38.955 ;
        RECT 117.365 37.345 119.035 38.435 ;
        RECT 119.205 38.145 119.515 39.155 ;
        RECT 119.685 38.535 119.855 38.985 ;
        RECT 120.025 38.705 120.415 38.985 ;
        RECT 120.600 38.655 120.845 38.985 ;
        RECT 119.685 38.365 120.475 38.535 ;
        RECT 119.205 37.515 119.645 38.145 ;
        RECT 119.820 37.345 120.135 38.195 ;
        RECT 120.305 37.685 120.475 38.365 ;
        RECT 120.645 37.855 120.845 38.655 ;
        RECT 121.045 37.855 121.295 38.985 ;
        RECT 121.510 38.655 121.915 38.985 ;
        RECT 122.085 38.485 122.255 39.155 ;
        RECT 122.430 39.130 122.885 39.895 ;
        RECT 123.160 39.515 124.460 39.725 ;
        RECT 124.715 39.535 125.045 39.895 ;
        RECT 124.290 39.365 124.460 39.515 ;
        RECT 125.215 39.395 125.475 39.725 ;
        RECT 123.360 38.905 123.580 39.305 ;
        RECT 122.425 38.705 122.915 38.905 ;
        RECT 123.105 38.695 123.580 38.905 ;
        RECT 123.825 38.905 124.035 39.305 ;
        RECT 124.290 39.240 125.045 39.365 ;
        RECT 124.290 39.195 125.135 39.240 ;
        RECT 124.865 39.075 125.135 39.195 ;
        RECT 123.825 38.695 124.155 38.905 ;
        RECT 124.325 38.635 124.735 38.940 ;
        RECT 121.485 38.315 122.255 38.485 ;
        RECT 122.430 38.465 123.605 38.525 ;
        RECT 124.965 38.500 125.135 39.075 ;
        RECT 124.935 38.465 125.135 38.500 ;
        RECT 122.430 38.355 125.135 38.465 ;
        RECT 121.485 37.685 121.735 38.315 ;
        RECT 120.305 37.515 121.735 37.685 ;
        RECT 121.915 37.345 122.245 38.145 ;
        RECT 122.430 37.735 122.685 38.355 ;
        RECT 123.275 38.295 125.075 38.355 ;
        RECT 123.275 38.265 123.605 38.295 ;
        RECT 125.305 38.195 125.475 39.395 ;
        RECT 125.650 39.130 126.105 39.895 ;
        RECT 126.380 39.515 127.680 39.725 ;
        RECT 127.935 39.535 128.265 39.895 ;
        RECT 127.510 39.365 127.680 39.515 ;
        RECT 128.435 39.395 128.695 39.725 ;
        RECT 126.580 38.905 126.800 39.305 ;
        RECT 125.645 38.705 126.135 38.905 ;
        RECT 126.325 38.695 126.800 38.905 ;
        RECT 127.045 38.905 127.255 39.305 ;
        RECT 127.510 39.240 128.265 39.365 ;
        RECT 127.510 39.195 128.355 39.240 ;
        RECT 128.085 39.075 128.355 39.195 ;
        RECT 127.045 38.695 127.375 38.905 ;
        RECT 127.545 38.635 127.955 38.940 ;
        RECT 122.935 38.095 123.120 38.185 ;
        RECT 123.710 38.095 124.545 38.105 ;
        RECT 122.935 37.895 124.545 38.095 ;
        RECT 122.935 37.855 123.165 37.895 ;
        RECT 122.430 37.515 122.765 37.735 ;
        RECT 123.770 37.345 124.125 37.725 ;
        RECT 124.295 37.515 124.545 37.895 ;
        RECT 124.795 37.345 125.045 38.125 ;
        RECT 125.215 37.515 125.475 38.195 ;
        RECT 125.650 38.465 126.825 38.525 ;
        RECT 128.185 38.500 128.355 39.075 ;
        RECT 128.155 38.465 128.355 38.500 ;
        RECT 125.650 38.355 128.355 38.465 ;
        RECT 125.650 37.735 125.905 38.355 ;
        RECT 126.495 38.295 128.295 38.355 ;
        RECT 126.495 38.265 126.825 38.295 ;
        RECT 128.525 38.195 128.695 39.395 ;
        RECT 128.875 39.245 129.205 39.710 ;
        RECT 129.375 39.425 129.545 39.895 ;
        RECT 129.720 39.495 130.050 39.725 ;
        RECT 129.800 39.245 129.970 39.495 ;
        RECT 130.255 39.335 130.425 39.725 ;
        RECT 128.875 39.075 129.970 39.245 ;
        RECT 130.185 39.155 130.425 39.335 ;
        RECT 130.770 39.325 130.960 39.485 ;
        RECT 130.650 39.155 130.960 39.325 ;
        RECT 131.180 39.155 131.455 39.895 ;
        RECT 128.865 38.695 129.345 38.905 ;
        RECT 129.515 38.695 130.015 38.905 ;
        RECT 130.185 38.525 130.355 39.155 ;
        RECT 130.650 38.985 130.820 39.155 ;
        RECT 131.685 39.075 131.895 39.895 ;
        RECT 132.065 39.095 132.395 39.725 ;
        RECT 126.155 38.095 126.340 38.185 ;
        RECT 126.930 38.095 127.765 38.105 ;
        RECT 126.155 37.895 127.765 38.095 ;
        RECT 126.155 37.855 126.385 37.895 ;
        RECT 125.650 37.515 125.985 37.735 ;
        RECT 126.990 37.345 127.345 37.725 ;
        RECT 127.515 37.515 127.765 37.895 ;
        RECT 128.015 37.345 128.265 38.125 ;
        RECT 128.435 37.515 128.695 38.195 ;
        RECT 128.895 37.345 129.270 38.445 ;
        RECT 129.745 38.355 130.355 38.525 ;
        RECT 130.525 38.445 130.820 38.985 ;
        RECT 131.005 38.635 131.455 38.985 ;
        RECT 129.745 37.515 130.070 38.355 ;
        RECT 130.525 38.275 131.015 38.445 ;
        RECT 130.240 37.345 130.570 38.105 ;
        RECT 130.740 37.770 131.015 38.275 ;
        RECT 131.185 37.535 131.455 38.635 ;
        RECT 132.065 38.495 132.315 39.095 ;
        RECT 132.565 39.075 132.795 39.895 ;
        RECT 133.005 39.125 135.595 39.895 ;
        RECT 136.230 39.435 136.485 39.895 ;
        RECT 136.660 39.265 136.990 39.665 ;
        RECT 132.485 38.655 132.815 38.905 ;
        RECT 133.005 38.605 134.215 39.125 ;
        RECT 136.290 39.095 136.990 39.265 ;
        RECT 137.160 39.115 137.360 39.895 ;
        RECT 138.115 39.515 138.445 39.895 ;
        RECT 137.595 39.155 138.005 39.325 ;
        RECT 131.685 37.345 131.895 38.485 ;
        RECT 132.065 37.515 132.395 38.495 ;
        RECT 132.565 37.345 132.795 38.485 ;
        RECT 134.385 38.435 135.595 38.955 ;
        RECT 133.005 37.345 135.595 38.435 ;
        RECT 136.290 38.145 136.520 39.095 ;
        RECT 137.835 38.985 138.005 39.155 ;
        RECT 138.485 39.155 138.880 39.345 ;
        RECT 139.375 39.155 139.705 39.895 ;
        RECT 139.915 39.165 140.215 39.895 ;
        RECT 137.470 38.945 137.665 38.985 ;
        RECT 136.710 38.485 137.040 38.905 ;
        RECT 137.210 38.655 137.665 38.945 ;
        RECT 137.835 38.655 138.315 38.985 ;
        RECT 136.710 38.315 137.425 38.485 ;
        RECT 137.835 38.425 138.005 38.655 ;
        RECT 138.485 38.475 138.655 39.155 ;
        RECT 140.395 38.985 140.625 39.605 ;
        RECT 140.825 39.335 141.050 39.715 ;
        RECT 141.220 39.505 141.550 39.895 ;
        RECT 140.825 39.155 141.155 39.335 ;
        RECT 136.290 37.975 136.990 38.145 ;
        RECT 136.230 37.345 136.565 37.725 ;
        RECT 136.735 37.555 136.990 37.975 ;
        RECT 137.255 38.085 137.425 38.315 ;
        RECT 137.595 38.255 138.005 38.425 ;
        RECT 138.195 38.305 138.655 38.475 ;
        RECT 138.825 38.365 139.240 38.985 ;
        RECT 139.410 38.365 139.700 38.985 ;
        RECT 139.920 38.655 140.215 38.985 ;
        RECT 140.395 38.655 140.810 38.985 ;
        RECT 140.980 38.485 141.155 39.155 ;
        RECT 141.325 38.655 141.565 39.305 ;
        RECT 142.665 39.170 142.955 39.895 ;
        RECT 143.175 39.505 143.505 39.895 ;
        RECT 143.675 39.325 143.845 39.645 ;
        RECT 144.015 39.505 144.345 39.895 ;
        RECT 144.760 39.495 145.715 39.665 ;
        RECT 143.125 39.155 145.375 39.325 ;
        RECT 138.195 38.085 138.365 38.305 ;
        RECT 137.255 37.875 138.365 38.085 ;
        RECT 137.180 37.345 137.510 37.705 ;
        RECT 138.115 37.515 138.365 37.875 ;
        RECT 138.535 37.965 139.705 38.135 ;
        RECT 138.535 37.515 138.865 37.965 ;
        RECT 139.035 37.345 139.205 37.795 ;
        RECT 139.375 37.515 139.705 37.965 ;
        RECT 139.915 38.125 140.810 38.455 ;
        RECT 140.980 38.295 141.565 38.485 ;
        RECT 139.915 37.955 141.120 38.125 ;
        RECT 139.915 37.525 140.245 37.955 ;
        RECT 140.425 37.345 140.620 37.785 ;
        RECT 140.790 37.525 141.120 37.955 ;
        RECT 141.290 37.525 141.565 38.295 ;
        RECT 142.665 37.345 142.955 38.510 ;
        RECT 143.125 38.195 143.295 39.155 ;
        RECT 143.465 38.535 143.710 38.985 ;
        RECT 143.880 38.705 144.430 38.905 ;
        RECT 144.600 38.735 144.975 38.905 ;
        RECT 144.600 38.535 144.770 38.735 ;
        RECT 145.145 38.655 145.375 39.155 ;
        RECT 143.465 38.365 144.770 38.535 ;
        RECT 145.545 38.615 145.715 39.495 ;
        RECT 145.885 39.060 146.175 39.895 ;
        RECT 147.265 39.155 147.650 39.725 ;
        RECT 147.820 39.435 148.145 39.895 ;
        RECT 148.665 39.265 148.945 39.725 ;
        RECT 145.545 38.445 146.175 38.615 ;
        RECT 143.125 37.515 143.505 38.195 ;
        RECT 144.095 37.345 144.265 38.195 ;
        RECT 144.435 38.025 145.675 38.195 ;
        RECT 144.435 37.515 144.765 38.025 ;
        RECT 144.935 37.345 145.105 37.855 ;
        RECT 145.275 37.515 145.675 38.025 ;
        RECT 145.855 37.515 146.175 38.445 ;
        RECT 147.265 38.485 147.545 39.155 ;
        RECT 147.820 39.095 148.945 39.265 ;
        RECT 147.820 38.985 148.270 39.095 ;
        RECT 147.715 38.655 148.270 38.985 ;
        RECT 149.135 38.925 149.535 39.725 ;
        RECT 149.935 39.435 150.205 39.895 ;
        RECT 150.375 39.265 150.660 39.725 ;
        RECT 147.265 37.515 147.650 38.485 ;
        RECT 147.820 38.195 148.270 38.655 ;
        RECT 148.440 38.365 149.535 38.925 ;
        RECT 147.820 37.975 148.945 38.195 ;
        RECT 147.820 37.345 148.145 37.805 ;
        RECT 148.665 37.515 148.945 37.975 ;
        RECT 149.135 37.515 149.535 38.365 ;
        RECT 149.705 39.095 150.660 39.265 ;
        RECT 150.945 39.145 152.155 39.895 ;
        RECT 149.705 38.195 149.915 39.095 ;
        RECT 150.085 38.365 150.775 38.925 ;
        RECT 150.945 38.435 151.465 38.975 ;
        RECT 151.635 38.605 152.155 39.145 ;
        RECT 149.705 37.975 150.660 38.195 ;
        RECT 149.935 37.345 150.205 37.805 ;
        RECT 150.375 37.515 150.660 37.975 ;
        RECT 150.945 37.345 152.155 38.435 ;
        RECT 91.060 37.175 152.240 37.345 ;
        RECT 91.145 36.085 92.355 37.175 ;
        RECT 91.145 35.375 91.665 35.915 ;
        RECT 91.835 35.545 92.355 36.085 ;
        RECT 92.530 36.035 92.785 37.175 ;
        RECT 92.980 36.625 94.175 36.955 ;
        RECT 93.035 35.865 93.205 36.425 ;
        RECT 93.430 36.205 93.850 36.455 ;
        RECT 94.355 36.375 94.635 37.175 ;
        RECT 93.430 36.035 94.675 36.205 ;
        RECT 94.845 36.035 95.115 37.005 ;
        RECT 95.285 36.665 95.545 37.175 ;
        RECT 94.505 35.865 94.675 36.035 ;
        RECT 92.530 35.615 92.865 35.865 ;
        RECT 93.035 35.535 93.775 35.865 ;
        RECT 94.505 35.535 94.735 35.865 ;
        RECT 93.035 35.445 93.285 35.535 ;
        RECT 6.025 33.760 6.380 34.100 ;
        RECT 6.030 31.940 6.380 33.760 ;
        RECT 59.055 32.505 59.405 34.665 ;
        RECT 91.145 34.625 92.355 35.375 ;
        RECT 92.550 35.275 93.285 35.445 ;
        RECT 94.505 35.365 94.675 35.535 ;
        RECT 92.550 34.805 92.860 35.275 ;
        RECT 93.935 35.195 94.675 35.365 ;
        RECT 94.945 35.300 95.115 36.035 ;
        RECT 95.285 35.615 95.625 36.495 ;
        RECT 95.795 35.785 95.965 37.005 ;
        RECT 96.205 36.670 96.820 37.175 ;
        RECT 96.205 36.135 96.455 36.500 ;
        RECT 96.625 36.495 96.820 36.670 ;
        RECT 96.990 36.665 97.465 37.005 ;
        RECT 97.635 36.630 97.850 37.175 ;
        RECT 96.625 36.305 96.955 36.495 ;
        RECT 97.175 36.135 97.890 36.430 ;
        RECT 98.060 36.305 98.335 37.005 ;
        RECT 98.505 36.375 98.830 37.175 ;
        RECT 96.205 35.965 97.995 36.135 ;
        RECT 95.795 35.535 96.590 35.785 ;
        RECT 95.795 35.445 96.045 35.535 ;
        RECT 93.030 34.625 93.765 35.105 ;
        RECT 93.935 34.845 94.105 35.195 ;
        RECT 94.275 34.625 94.655 35.025 ;
        RECT 94.845 34.955 95.115 35.300 ;
        RECT 95.285 34.625 95.545 35.445 ;
        RECT 95.715 35.025 96.045 35.445 ;
        RECT 96.760 35.110 97.015 35.965 ;
        RECT 96.225 34.845 97.015 35.110 ;
        RECT 97.185 35.265 97.595 35.785 ;
        RECT 97.765 35.535 97.995 35.965 ;
        RECT 98.165 35.275 98.335 36.305 ;
        RECT 98.525 35.615 98.855 36.200 ;
        RECT 99.025 35.865 99.210 36.955 ;
        RECT 99.380 36.205 99.630 37.005 ;
        RECT 99.800 36.375 100.540 37.175 ;
        RECT 100.725 36.205 101.055 37.005 ;
        RECT 101.225 36.375 102.035 37.175 ;
        RECT 99.380 36.035 101.865 36.205 ;
        RECT 101.695 35.865 101.865 36.035 ;
        RECT 99.025 35.615 99.510 35.865 ;
        RECT 99.855 35.535 100.115 35.865 ;
        RECT 97.185 34.845 97.385 35.265 ;
        RECT 97.575 34.625 97.905 35.085 ;
        RECT 98.075 34.795 98.335 35.275 ;
        RECT 98.505 35.245 99.690 35.415 ;
        RECT 98.505 34.795 98.770 35.245 ;
        RECT 98.940 34.625 99.230 35.075 ;
        RECT 99.400 34.795 99.690 35.245 ;
        RECT 99.870 34.930 100.115 35.535 ;
        RECT 100.365 34.930 100.635 35.865 ;
        RECT 100.815 35.615 101.295 35.865 ;
        RECT 100.815 34.930 101.025 35.615 ;
        RECT 101.695 35.535 102.035 35.865 ;
        RECT 101.695 35.445 101.865 35.535 ;
        RECT 101.195 35.275 101.865 35.445 ;
        RECT 101.195 34.795 101.535 35.275 ;
        RECT 101.715 34.625 102.025 35.105 ;
        RECT 102.205 34.795 102.465 37.005 ;
        RECT 102.685 36.035 102.915 37.175 ;
        RECT 103.085 36.025 103.415 37.005 ;
        RECT 103.585 36.035 103.795 37.175 ;
        RECT 102.665 35.615 102.995 35.865 ;
        RECT 102.685 34.625 102.915 35.445 ;
        RECT 103.165 35.425 103.415 36.025 ;
        RECT 104.025 36.010 104.315 37.175 ;
        RECT 104.640 36.165 104.940 37.005 ;
        RECT 105.135 36.335 105.385 37.175 ;
        RECT 105.975 36.585 106.780 37.005 ;
        RECT 105.555 36.415 107.120 36.585 ;
        RECT 105.555 36.165 105.725 36.415 ;
        RECT 104.640 35.995 105.725 36.165 ;
        RECT 104.485 35.535 104.815 35.825 ;
        RECT 103.085 34.795 103.415 35.425 ;
        RECT 103.585 34.625 103.795 35.445 ;
        RECT 104.985 35.365 105.155 35.995 ;
        RECT 105.895 35.865 106.215 36.245 ;
        RECT 106.405 36.155 106.780 36.245 ;
        RECT 106.385 35.985 106.780 36.155 ;
        RECT 106.950 36.165 107.120 36.415 ;
        RECT 107.290 36.335 107.620 37.175 ;
        RECT 107.790 36.415 108.455 37.005 ;
        RECT 106.950 35.995 107.870 36.165 ;
        RECT 105.325 35.615 105.655 35.825 ;
        RECT 105.835 35.615 106.215 35.865 ;
        RECT 106.405 35.825 106.780 35.985 ;
        RECT 107.700 35.825 107.870 35.995 ;
        RECT 106.405 35.615 106.890 35.825 ;
        RECT 107.080 35.615 107.530 35.825 ;
        RECT 107.700 35.615 108.035 35.825 ;
        RECT 108.205 35.445 108.455 36.415 ;
        RECT 109.700 36.165 110.000 37.005 ;
        RECT 110.195 36.335 110.445 37.175 ;
        RECT 111.035 36.585 111.840 37.005 ;
        RECT 110.615 36.415 112.180 36.585 ;
        RECT 110.615 36.165 110.785 36.415 ;
        RECT 109.700 35.995 110.785 36.165 ;
        RECT 109.545 35.535 109.875 35.825 ;
        RECT 104.025 34.625 104.315 35.350 ;
        RECT 104.645 35.185 105.155 35.365 ;
        RECT 105.560 35.275 107.260 35.445 ;
        RECT 105.560 35.185 105.945 35.275 ;
        RECT 104.645 34.795 104.975 35.185 ;
        RECT 105.145 34.845 106.330 35.015 ;
        RECT 106.590 34.625 106.760 35.095 ;
        RECT 106.930 34.810 107.260 35.275 ;
        RECT 107.430 34.625 107.600 35.445 ;
        RECT 107.770 34.805 108.455 35.445 ;
        RECT 110.045 35.365 110.215 35.995 ;
        RECT 110.955 35.865 111.275 36.245 ;
        RECT 111.465 36.155 111.840 36.245 ;
        RECT 111.445 35.985 111.840 36.155 ;
        RECT 112.010 36.165 112.180 36.415 ;
        RECT 112.350 36.335 112.680 37.175 ;
        RECT 112.850 36.415 113.515 37.005 ;
        RECT 112.010 35.995 112.930 36.165 ;
        RECT 110.385 35.615 110.715 35.825 ;
        RECT 110.895 35.615 111.275 35.865 ;
        RECT 111.465 35.825 111.840 35.985 ;
        RECT 112.760 35.825 112.930 35.995 ;
        RECT 111.465 35.615 111.950 35.825 ;
        RECT 112.140 35.615 112.590 35.825 ;
        RECT 112.760 35.615 113.095 35.825 ;
        RECT 113.265 35.445 113.515 36.415 ;
        RECT 113.745 36.035 113.955 37.175 ;
        RECT 114.125 36.025 114.455 37.005 ;
        RECT 114.625 36.035 114.855 37.175 ;
        RECT 109.705 35.185 110.215 35.365 ;
        RECT 110.620 35.275 112.320 35.445 ;
        RECT 110.620 35.185 111.005 35.275 ;
        RECT 109.705 34.795 110.035 35.185 ;
        RECT 110.205 34.845 111.390 35.015 ;
        RECT 111.650 34.625 111.820 35.095 ;
        RECT 111.990 34.810 112.320 35.275 ;
        RECT 112.490 34.625 112.660 35.445 ;
        RECT 112.830 34.805 113.515 35.445 ;
        RECT 113.745 34.625 113.955 35.445 ;
        RECT 114.125 35.425 114.375 36.025 ;
        RECT 114.545 35.615 114.875 35.865 ;
        RECT 114.125 34.795 114.455 35.425 ;
        RECT 114.625 34.625 114.855 35.445 ;
        RECT 115.065 34.905 115.345 37.005 ;
        RECT 115.535 36.415 116.320 37.175 ;
        RECT 116.715 36.345 117.100 37.005 ;
        RECT 116.715 36.245 117.125 36.345 ;
        RECT 115.515 36.035 117.125 36.245 ;
        RECT 117.425 36.155 117.625 36.945 ;
        RECT 115.515 35.435 115.790 36.035 ;
        RECT 117.295 35.985 117.625 36.155 ;
        RECT 117.795 35.995 118.115 37.175 ;
        RECT 118.285 36.085 119.955 37.175 ;
        RECT 120.130 36.665 121.785 36.955 ;
        RECT 117.295 35.865 117.475 35.985 ;
        RECT 115.960 35.615 116.315 35.865 ;
        RECT 116.510 35.815 116.975 35.865 ;
        RECT 116.505 35.645 116.975 35.815 ;
        RECT 116.510 35.615 116.975 35.645 ;
        RECT 117.145 35.615 117.475 35.865 ;
        RECT 117.650 35.615 118.115 35.815 ;
        RECT 115.515 35.255 116.765 35.435 ;
        RECT 116.400 35.185 116.765 35.255 ;
        RECT 116.935 35.235 118.115 35.405 ;
        RECT 115.575 34.625 115.745 35.085 ;
        RECT 116.935 35.015 117.265 35.235 ;
        RECT 116.015 34.835 117.265 35.015 ;
        RECT 117.435 34.625 117.605 35.065 ;
        RECT 117.775 34.820 118.115 35.235 ;
        RECT 118.285 35.395 119.035 35.915 ;
        RECT 119.205 35.565 119.955 36.085 ;
        RECT 120.130 36.325 121.720 36.495 ;
        RECT 121.955 36.375 122.235 37.175 ;
        RECT 120.130 36.035 120.450 36.325 ;
        RECT 121.550 36.205 121.720 36.325 ;
        RECT 118.285 34.625 119.955 35.395 ;
        RECT 120.130 35.295 120.480 35.865 ;
        RECT 120.650 35.535 121.360 36.155 ;
        RECT 121.550 36.035 122.275 36.205 ;
        RECT 122.445 36.035 122.715 37.005 ;
        RECT 122.105 35.865 122.275 36.035 ;
        RECT 121.530 35.535 121.935 35.865 ;
        RECT 122.105 35.535 122.375 35.865 ;
        RECT 122.105 35.365 122.275 35.535 ;
        RECT 120.665 35.195 122.275 35.365 ;
        RECT 122.545 35.300 122.715 36.035 ;
        RECT 120.135 34.625 120.465 35.125 ;
        RECT 120.665 34.845 120.835 35.195 ;
        RECT 121.035 34.625 121.365 35.025 ;
        RECT 121.535 34.845 121.705 35.195 ;
        RECT 121.875 34.625 122.255 35.025 ;
        RECT 122.445 34.955 122.715 35.300 ;
        RECT 122.885 36.335 123.145 37.005 ;
        RECT 123.315 36.775 123.645 37.175 ;
        RECT 124.515 36.775 124.915 37.175 ;
        RECT 125.205 36.595 125.535 36.830 ;
        RECT 123.455 36.425 125.535 36.595 ;
        RECT 122.885 35.365 123.060 36.335 ;
        RECT 123.455 36.155 123.625 36.425 ;
        RECT 123.230 35.985 123.625 36.155 ;
        RECT 123.795 36.035 124.810 36.255 ;
        RECT 123.230 35.535 123.400 35.985 ;
        RECT 124.535 35.895 124.810 36.035 ;
        RECT 124.980 36.035 125.535 36.425 ;
        RECT 123.570 35.615 124.020 35.815 ;
        RECT 124.190 35.445 124.365 35.640 ;
        RECT 122.885 34.795 123.225 35.365 ;
        RECT 123.420 34.625 123.590 35.290 ;
        RECT 123.870 35.275 124.365 35.445 ;
        RECT 123.870 35.135 124.090 35.275 ;
        RECT 123.865 34.965 124.090 35.135 ;
        RECT 124.535 35.105 124.705 35.895 ;
        RECT 124.980 35.785 125.150 36.035 ;
        RECT 125.705 35.865 125.880 36.965 ;
        RECT 126.050 36.355 126.395 37.175 ;
        RECT 126.565 36.325 126.825 37.005 ;
        RECT 126.995 36.395 127.245 37.175 ;
        RECT 127.495 36.625 127.745 37.005 ;
        RECT 127.915 36.795 128.270 37.175 ;
        RECT 129.275 36.785 129.610 37.005 ;
        RECT 128.875 36.625 129.105 36.665 ;
        RECT 127.495 36.425 129.105 36.625 ;
        RECT 127.495 36.415 128.330 36.425 ;
        RECT 128.920 36.335 129.105 36.425 ;
        RECT 124.955 35.615 125.150 35.785 ;
        RECT 125.320 35.615 125.880 35.865 ;
        RECT 126.050 35.615 126.395 36.185 ;
        RECT 124.955 35.230 125.125 35.615 ;
        RECT 123.870 34.920 124.090 34.965 ;
        RECT 124.260 34.935 124.705 35.105 ;
        RECT 124.875 34.860 125.125 35.230 ;
        RECT 125.295 35.265 126.395 35.445 ;
        RECT 125.295 34.860 125.545 35.265 ;
        RECT 125.715 34.625 125.885 35.095 ;
        RECT 126.055 34.860 126.395 35.265 ;
        RECT 126.565 35.135 126.735 36.325 ;
        RECT 128.435 36.225 128.765 36.255 ;
        RECT 126.965 36.165 128.765 36.225 ;
        RECT 129.355 36.165 129.610 36.785 ;
        RECT 126.905 36.055 129.610 36.165 ;
        RECT 126.905 36.020 127.105 36.055 ;
        RECT 126.905 35.445 127.075 36.020 ;
        RECT 128.435 35.995 129.610 36.055 ;
        RECT 129.785 36.010 130.075 37.175 ;
        RECT 127.305 35.580 127.715 35.885 ;
        RECT 127.885 35.615 128.215 35.825 ;
        RECT 126.905 35.325 127.175 35.445 ;
        RECT 126.905 35.280 127.750 35.325 ;
        RECT 126.995 35.155 127.750 35.280 ;
        RECT 128.005 35.215 128.215 35.615 ;
        RECT 128.460 35.615 128.935 35.825 ;
        RECT 129.125 35.615 129.615 35.815 ;
        RECT 128.460 35.215 128.680 35.615 ;
        RECT 126.565 35.125 126.795 35.135 ;
        RECT 126.565 34.795 126.825 35.125 ;
        RECT 127.580 35.005 127.750 35.155 ;
        RECT 126.995 34.625 127.325 34.985 ;
        RECT 127.580 34.795 128.880 35.005 ;
        RECT 129.155 34.625 129.610 35.390 ;
        RECT 129.785 34.625 130.075 35.350 ;
        RECT 130.245 34.905 130.525 37.005 ;
        RECT 130.715 36.415 131.500 37.175 ;
        RECT 131.895 36.345 132.280 37.005 ;
        RECT 131.895 36.245 132.305 36.345 ;
        RECT 130.695 36.035 132.305 36.245 ;
        RECT 132.605 36.155 132.805 36.945 ;
        RECT 130.695 35.435 130.970 36.035 ;
        RECT 132.475 35.985 132.805 36.155 ;
        RECT 132.975 35.995 133.295 37.175 ;
        RECT 133.555 36.165 133.725 37.005 ;
        RECT 133.895 36.835 135.065 37.005 ;
        RECT 133.895 36.335 134.225 36.835 ;
        RECT 134.735 36.795 135.065 36.835 ;
        RECT 135.255 36.755 135.610 37.175 ;
        RECT 134.395 36.575 134.625 36.665 ;
        RECT 135.780 36.575 136.030 37.005 ;
        RECT 134.395 36.335 136.030 36.575 ;
        RECT 136.200 36.415 136.530 37.175 ;
        RECT 136.700 36.335 136.955 37.005 ;
        RECT 133.555 35.995 136.615 36.165 ;
        RECT 132.475 35.865 132.655 35.985 ;
        RECT 131.140 35.615 131.495 35.865 ;
        RECT 131.690 35.815 132.155 35.865 ;
        RECT 131.685 35.645 132.155 35.815 ;
        RECT 131.690 35.615 132.155 35.645 ;
        RECT 132.325 35.615 132.655 35.865 ;
        RECT 132.830 35.615 133.295 35.815 ;
        RECT 133.470 35.615 133.820 35.825 ;
        RECT 133.990 35.615 134.435 35.815 ;
        RECT 134.605 35.615 135.080 35.815 ;
        RECT 130.695 35.255 131.945 35.435 ;
        RECT 131.580 35.185 131.945 35.255 ;
        RECT 132.115 35.235 133.295 35.405 ;
        RECT 130.755 34.625 130.925 35.085 ;
        RECT 132.115 35.015 132.445 35.235 ;
        RECT 131.195 34.835 132.445 35.015 ;
        RECT 132.615 34.625 132.785 35.065 ;
        RECT 132.955 34.820 133.295 35.235 ;
        RECT 133.555 35.275 134.620 35.445 ;
        RECT 133.555 34.795 133.725 35.275 ;
        RECT 133.895 34.625 134.225 35.105 ;
        RECT 134.450 35.045 134.620 35.275 ;
        RECT 134.800 35.215 135.080 35.615 ;
        RECT 135.350 35.615 135.680 35.815 ;
        RECT 135.850 35.615 136.215 35.815 ;
        RECT 135.350 35.215 135.635 35.615 ;
        RECT 136.445 35.445 136.615 35.995 ;
        RECT 135.815 35.275 136.615 35.445 ;
        RECT 135.815 35.045 135.985 35.275 ;
        RECT 136.785 35.205 136.955 36.335 ;
        RECT 137.615 36.035 137.945 37.175 ;
        RECT 138.475 36.205 138.805 36.990 ;
        RECT 138.125 36.035 138.805 36.205 ;
        RECT 139.945 36.035 140.175 37.175 ;
        RECT 137.605 35.615 137.955 35.865 ;
        RECT 138.125 35.435 138.295 36.035 ;
        RECT 140.345 36.025 140.675 37.005 ;
        RECT 140.845 36.035 141.055 37.175 ;
        RECT 141.290 36.505 141.545 37.005 ;
        RECT 141.715 36.675 142.045 37.175 ;
        RECT 141.290 36.335 142.040 36.505 ;
        RECT 138.465 35.615 138.815 35.865 ;
        RECT 139.925 35.615 140.255 35.865 ;
        RECT 136.770 35.125 136.955 35.205 ;
        RECT 134.450 34.795 135.985 35.045 ;
        RECT 136.155 34.625 136.485 35.105 ;
        RECT 136.700 34.795 136.955 35.125 ;
        RECT 137.615 34.625 137.885 35.435 ;
        RECT 138.055 34.795 138.385 35.435 ;
        RECT 138.555 34.625 138.795 35.435 ;
        RECT 139.945 34.625 140.175 35.445 ;
        RECT 140.425 35.425 140.675 36.025 ;
        RECT 141.290 35.515 141.640 36.165 ;
        RECT 140.345 34.795 140.675 35.425 ;
        RECT 140.845 34.625 141.055 35.445 ;
        RECT 141.810 35.345 142.040 36.335 ;
        RECT 141.290 35.175 142.040 35.345 ;
        RECT 141.290 34.885 141.545 35.175 ;
        RECT 141.715 34.625 142.045 35.005 ;
        RECT 142.215 34.885 142.385 37.005 ;
        RECT 142.555 36.205 142.880 36.990 ;
        RECT 143.050 36.715 143.300 37.175 ;
        RECT 143.470 36.675 143.720 37.005 ;
        RECT 143.935 36.675 144.615 37.005 ;
        RECT 143.470 36.545 143.640 36.675 ;
        RECT 143.245 36.375 143.640 36.545 ;
        RECT 142.615 35.155 143.075 36.205 ;
        RECT 143.245 35.015 143.415 36.375 ;
        RECT 143.810 36.115 144.275 36.505 ;
        RECT 143.585 35.305 143.935 35.925 ;
        RECT 144.105 35.525 144.275 36.115 ;
        RECT 144.445 35.895 144.615 36.675 ;
        RECT 144.785 36.575 144.955 36.915 ;
        RECT 145.190 36.745 145.520 37.175 ;
        RECT 145.690 36.575 145.860 36.915 ;
        RECT 146.155 36.715 146.525 37.175 ;
        RECT 144.785 36.405 145.860 36.575 ;
        RECT 146.695 36.545 146.865 37.005 ;
        RECT 147.100 36.665 147.970 37.005 ;
        RECT 148.140 36.715 148.390 37.175 ;
        RECT 146.305 36.375 146.865 36.545 ;
        RECT 146.305 36.235 146.475 36.375 ;
        RECT 144.975 36.065 146.475 36.235 ;
        RECT 147.170 36.205 147.630 36.495 ;
        RECT 144.445 35.725 146.135 35.895 ;
        RECT 144.105 35.305 144.460 35.525 ;
        RECT 144.630 35.015 144.800 35.725 ;
        RECT 145.005 35.305 145.795 35.555 ;
        RECT 145.965 35.545 146.135 35.725 ;
        RECT 146.305 35.375 146.475 36.065 ;
        RECT 142.745 34.625 143.075 34.985 ;
        RECT 143.245 34.845 143.740 35.015 ;
        RECT 143.945 34.845 144.800 35.015 ;
        RECT 145.675 34.625 146.005 35.085 ;
        RECT 146.215 34.985 146.475 35.375 ;
        RECT 146.665 36.195 147.630 36.205 ;
        RECT 147.800 36.285 147.970 36.665 ;
        RECT 148.560 36.625 148.730 36.915 ;
        RECT 148.910 36.795 149.240 37.175 ;
        RECT 148.560 36.455 149.360 36.625 ;
        RECT 146.665 36.035 147.340 36.195 ;
        RECT 147.800 36.115 149.020 36.285 ;
        RECT 146.665 35.245 146.875 36.035 ;
        RECT 147.800 36.025 147.970 36.115 ;
        RECT 147.045 35.245 147.395 35.865 ;
        RECT 147.565 35.855 147.970 36.025 ;
        RECT 147.565 35.075 147.735 35.855 ;
        RECT 147.905 35.405 148.125 35.685 ;
        RECT 148.305 35.575 148.845 35.945 ;
        RECT 149.190 35.865 149.360 36.455 ;
        RECT 149.580 36.035 149.885 37.175 ;
        RECT 150.055 35.985 150.310 36.865 ;
        RECT 149.190 35.835 149.930 35.865 ;
        RECT 147.905 35.235 148.435 35.405 ;
        RECT 146.215 34.815 146.565 34.985 ;
        RECT 146.785 34.795 147.735 35.075 ;
        RECT 147.905 34.625 148.095 35.065 ;
        RECT 148.265 35.005 148.435 35.235 ;
        RECT 148.605 35.175 148.845 35.575 ;
        RECT 149.015 35.535 149.930 35.835 ;
        RECT 149.015 35.360 149.340 35.535 ;
        RECT 149.015 35.005 149.335 35.360 ;
        RECT 150.100 35.335 150.310 35.985 ;
        RECT 150.945 36.085 152.155 37.175 ;
        RECT 150.945 35.545 151.465 36.085 ;
        RECT 151.635 35.375 152.155 35.915 ;
        RECT 148.265 34.835 149.335 35.005 ;
        RECT 149.580 34.625 149.885 35.085 ;
        RECT 150.055 34.805 150.310 35.335 ;
        RECT 150.945 34.625 152.155 35.375 ;
        RECT 91.060 34.455 152.240 34.625 ;
        RECT 91.145 33.705 92.355 34.455 ;
        RECT 92.525 33.910 97.870 34.455 ;
        RECT 91.145 33.165 91.665 33.705 ;
        RECT 91.835 32.995 92.355 33.535 ;
        RECT 94.110 33.080 94.450 33.910 ;
        RECT 98.070 33.805 98.380 34.275 ;
        RECT 98.550 33.975 99.285 34.455 ;
        RECT 99.455 33.885 99.625 34.235 ;
        RECT 99.795 34.055 100.175 34.455 ;
        RECT 98.070 33.635 98.805 33.805 ;
        RECT 99.455 33.715 100.195 33.885 ;
        RECT 100.365 33.780 100.635 34.125 ;
        RECT 91.145 31.905 92.355 32.995 ;
        RECT 95.930 32.340 96.280 33.590 ;
        RECT 98.555 33.545 98.805 33.635 ;
        RECT 100.025 33.545 100.195 33.715 ;
        RECT 98.050 33.215 98.385 33.465 ;
        RECT 98.555 33.215 99.295 33.545 ;
        RECT 100.025 33.215 100.255 33.545 ;
        RECT 92.525 31.905 97.870 32.340 ;
        RECT 98.050 31.905 98.305 33.045 ;
        RECT 98.555 32.655 98.725 33.215 ;
        RECT 100.025 33.045 100.195 33.215 ;
        RECT 100.465 33.045 100.635 33.780 ;
        RECT 98.950 32.875 100.195 33.045 ;
        RECT 98.950 32.625 99.370 32.875 ;
        RECT 98.500 32.125 99.695 32.455 ;
        RECT 99.875 31.905 100.155 32.705 ;
        RECT 100.365 32.075 100.635 33.045 ;
        RECT 100.805 33.780 101.075 34.125 ;
        RECT 101.265 34.055 101.645 34.455 ;
        RECT 101.815 33.885 101.985 34.235 ;
        RECT 102.155 33.975 102.890 34.455 ;
        RECT 100.805 33.045 100.975 33.780 ;
        RECT 101.245 33.715 101.985 33.885 ;
        RECT 103.060 33.805 103.370 34.275 ;
        RECT 101.245 33.545 101.415 33.715 ;
        RECT 102.635 33.635 103.370 33.805 ;
        RECT 104.025 33.870 104.335 34.285 ;
        RECT 104.530 34.075 104.860 34.455 ;
        RECT 105.030 34.115 106.435 34.285 ;
        RECT 105.030 33.885 105.200 34.115 ;
        RECT 102.635 33.545 102.885 33.635 ;
        RECT 101.185 33.215 101.415 33.545 ;
        RECT 102.145 33.215 102.885 33.545 ;
        RECT 103.055 33.215 103.390 33.465 ;
        RECT 101.245 33.045 101.415 33.215 ;
        RECT 100.805 32.075 101.075 33.045 ;
        RECT 101.245 32.875 102.490 33.045 ;
        RECT 101.285 31.905 101.565 32.705 ;
        RECT 102.070 32.625 102.490 32.875 ;
        RECT 102.715 32.655 102.885 33.215 ;
        RECT 101.745 32.125 102.940 32.455 ;
        RECT 103.135 31.905 103.390 33.045 ;
        RECT 104.025 32.755 104.195 33.870 ;
        RECT 104.505 33.715 105.200 33.885 ;
        RECT 106.265 33.885 106.435 34.115 ;
        RECT 106.705 34.055 107.035 34.455 ;
        RECT 107.275 33.885 107.445 34.285 ;
        RECT 104.505 33.545 104.675 33.715 ;
        RECT 104.365 33.215 104.675 33.545 ;
        RECT 104.845 33.215 105.180 33.545 ;
        RECT 105.450 33.215 105.645 33.790 ;
        RECT 105.905 33.545 106.095 33.775 ;
        RECT 106.265 33.715 107.445 33.885 ;
        RECT 107.725 33.765 107.965 34.285 ;
        RECT 108.135 33.960 108.530 34.455 ;
        RECT 109.095 34.125 109.265 34.270 ;
        RECT 108.890 33.930 109.265 34.125 ;
        RECT 105.905 33.215 106.250 33.545 ;
        RECT 106.560 33.215 107.035 33.545 ;
        RECT 107.290 33.215 107.475 33.545 ;
        RECT 104.505 33.045 104.675 33.215 ;
        RECT 104.505 32.875 107.445 33.045 ;
        RECT 104.025 32.115 104.365 32.755 ;
        RECT 104.955 32.535 106.515 32.705 ;
        RECT 104.535 31.905 104.780 32.365 ;
        RECT 104.955 32.075 105.205 32.535 ;
        RECT 105.395 31.905 106.065 32.285 ;
        RECT 106.265 32.075 106.515 32.535 ;
        RECT 107.275 32.075 107.445 32.875 ;
        RECT 107.725 32.960 107.900 33.765 ;
        RECT 108.890 33.595 109.060 33.930 ;
        RECT 109.545 33.885 109.785 34.260 ;
        RECT 109.955 33.950 110.290 34.455 ;
        RECT 109.545 33.735 109.765 33.885 ;
        RECT 108.075 33.235 109.060 33.595 ;
        RECT 109.230 33.405 109.765 33.735 ;
        RECT 108.075 33.215 109.360 33.235 ;
        RECT 108.500 33.065 109.360 33.215 ;
        RECT 107.725 32.175 108.030 32.960 ;
        RECT 108.205 32.585 108.900 32.895 ;
        RECT 108.210 31.905 108.895 32.375 ;
        RECT 109.075 32.120 109.360 33.065 ;
        RECT 109.530 32.755 109.765 33.405 ;
        RECT 109.935 32.925 110.235 33.775 ;
        RECT 110.930 33.690 111.385 34.455 ;
        RECT 111.660 34.075 112.960 34.285 ;
        RECT 113.215 34.095 113.545 34.455 ;
        RECT 112.790 33.925 112.960 34.075 ;
        RECT 113.715 33.955 113.975 34.285 ;
        RECT 113.745 33.945 113.975 33.955 ;
        RECT 111.860 33.465 112.080 33.865 ;
        RECT 110.925 33.265 111.415 33.465 ;
        RECT 111.605 33.255 112.080 33.465 ;
        RECT 112.325 33.465 112.535 33.865 ;
        RECT 112.790 33.800 113.545 33.925 ;
        RECT 112.790 33.755 113.635 33.800 ;
        RECT 113.365 33.635 113.635 33.755 ;
        RECT 112.325 33.255 112.655 33.465 ;
        RECT 112.825 33.195 113.235 33.500 ;
        RECT 110.930 33.025 112.105 33.085 ;
        RECT 113.465 33.060 113.635 33.635 ;
        RECT 113.435 33.025 113.635 33.060 ;
        RECT 110.930 32.915 113.635 33.025 ;
        RECT 109.530 32.525 110.205 32.755 ;
        RECT 109.535 31.905 109.865 32.355 ;
        RECT 110.035 32.095 110.205 32.525 ;
        RECT 110.930 32.295 111.185 32.915 ;
        RECT 111.775 32.855 113.575 32.915 ;
        RECT 111.775 32.825 112.105 32.855 ;
        RECT 113.805 32.755 113.975 33.945 ;
        RECT 111.435 32.655 111.620 32.745 ;
        RECT 112.210 32.655 113.045 32.665 ;
        RECT 111.435 32.455 113.045 32.655 ;
        RECT 111.435 32.415 111.665 32.455 ;
        RECT 110.930 32.075 111.265 32.295 ;
        RECT 112.270 31.905 112.625 32.285 ;
        RECT 112.795 32.075 113.045 32.455 ;
        RECT 113.295 31.905 113.545 32.685 ;
        RECT 113.715 32.075 113.975 32.755 ;
        RECT 114.180 33.715 114.795 34.285 ;
        RECT 114.965 33.945 115.180 34.455 ;
        RECT 115.410 33.945 115.690 34.275 ;
        RECT 115.870 33.945 116.110 34.455 ;
        RECT 114.180 32.695 114.495 33.715 ;
        RECT 114.665 33.045 114.835 33.545 ;
        RECT 115.085 33.215 115.350 33.775 ;
        RECT 115.520 33.045 115.690 33.945 ;
        RECT 115.860 33.215 116.215 33.775 ;
        RECT 116.905 33.730 117.195 34.455 ;
        RECT 117.835 33.955 118.165 34.455 ;
        RECT 118.365 33.885 118.535 34.235 ;
        RECT 118.735 34.055 119.065 34.455 ;
        RECT 119.235 33.885 119.405 34.235 ;
        RECT 119.575 34.055 119.955 34.455 ;
        RECT 117.830 33.215 118.180 33.785 ;
        RECT 118.365 33.715 119.975 33.885 ;
        RECT 120.145 33.780 120.415 34.125 ;
        RECT 119.805 33.545 119.975 33.715 ;
        RECT 114.665 32.875 116.090 33.045 ;
        RECT 114.180 32.075 114.715 32.695 ;
        RECT 114.885 31.905 115.215 32.705 ;
        RECT 115.700 32.700 116.090 32.875 ;
        RECT 116.905 31.905 117.195 33.070 ;
        RECT 117.830 32.755 118.150 33.045 ;
        RECT 118.350 32.925 119.060 33.545 ;
        RECT 119.230 33.215 119.635 33.545 ;
        RECT 119.805 33.215 120.075 33.545 ;
        RECT 119.805 33.045 119.975 33.215 ;
        RECT 120.245 33.045 120.415 33.780 ;
        RECT 121.565 33.635 121.775 34.455 ;
        RECT 121.945 33.655 122.275 34.285 ;
        RECT 121.945 33.055 122.195 33.655 ;
        RECT 122.445 33.635 122.675 34.455 ;
        RECT 122.905 33.725 123.195 34.455 ;
        RECT 122.365 33.215 122.695 33.465 ;
        RECT 122.895 33.215 123.195 33.545 ;
        RECT 123.375 33.525 123.605 34.165 ;
        RECT 123.785 33.905 124.095 34.275 ;
        RECT 124.275 34.085 124.945 34.455 ;
        RECT 123.785 33.705 125.015 33.905 ;
        RECT 123.375 33.215 123.900 33.525 ;
        RECT 124.080 33.215 124.545 33.525 ;
        RECT 119.250 32.875 119.975 33.045 ;
        RECT 119.250 32.755 119.420 32.875 ;
        RECT 117.830 32.585 119.420 32.755 ;
        RECT 117.830 32.125 119.485 32.415 ;
        RECT 119.655 31.905 119.935 32.705 ;
        RECT 120.145 32.075 120.415 33.045 ;
        RECT 121.565 31.905 121.775 33.045 ;
        RECT 121.945 32.075 122.275 33.055 ;
        RECT 122.445 31.905 122.675 33.045 ;
        RECT 124.725 33.035 125.015 33.705 ;
        RECT 122.905 32.795 124.065 33.035 ;
        RECT 122.905 32.085 123.165 32.795 ;
        RECT 123.335 31.905 123.665 32.615 ;
        RECT 123.835 32.085 124.065 32.795 ;
        RECT 124.245 32.815 125.015 33.035 ;
        RECT 124.245 32.085 124.515 32.815 ;
        RECT 124.695 31.905 125.035 32.635 ;
        RECT 125.205 32.085 125.465 34.275 ;
        RECT 126.570 33.690 127.025 34.455 ;
        RECT 127.300 34.075 128.600 34.285 ;
        RECT 128.855 34.095 129.185 34.455 ;
        RECT 128.430 33.925 128.600 34.075 ;
        RECT 129.355 33.955 129.615 34.285 ;
        RECT 129.385 33.945 129.615 33.955 ;
        RECT 127.500 33.465 127.720 33.865 ;
        RECT 126.565 33.265 127.055 33.465 ;
        RECT 127.245 33.255 127.720 33.465 ;
        RECT 127.965 33.465 128.175 33.865 ;
        RECT 128.430 33.800 129.185 33.925 ;
        RECT 128.430 33.755 129.275 33.800 ;
        RECT 129.005 33.635 129.275 33.755 ;
        RECT 127.965 33.255 128.295 33.465 ;
        RECT 128.465 33.195 128.875 33.500 ;
        RECT 126.570 33.025 127.745 33.085 ;
        RECT 129.105 33.060 129.275 33.635 ;
        RECT 129.075 33.025 129.275 33.060 ;
        RECT 126.570 32.915 129.275 33.025 ;
        RECT 126.570 32.295 126.825 32.915 ;
        RECT 127.415 32.855 129.215 32.915 ;
        RECT 127.415 32.825 127.745 32.855 ;
        RECT 129.445 32.755 129.615 33.945 ;
        RECT 129.785 33.705 130.995 34.455 ;
        RECT 131.165 33.845 131.505 34.260 ;
        RECT 131.675 34.015 131.845 34.455 ;
        RECT 132.015 34.065 133.265 34.245 ;
        RECT 132.015 33.845 132.345 34.065 ;
        RECT 133.535 33.995 133.705 34.455 ;
        RECT 129.785 33.165 130.305 33.705 ;
        RECT 131.165 33.675 132.345 33.845 ;
        RECT 132.515 33.825 132.880 33.895 ;
        RECT 132.515 33.645 133.765 33.825 ;
        RECT 130.475 32.995 130.995 33.535 ;
        RECT 131.165 33.265 131.630 33.465 ;
        RECT 131.805 33.215 132.135 33.465 ;
        RECT 132.305 33.435 132.770 33.465 ;
        RECT 132.305 33.265 132.775 33.435 ;
        RECT 132.305 33.215 132.770 33.265 ;
        RECT 132.965 33.215 133.320 33.465 ;
        RECT 131.805 33.095 131.985 33.215 ;
        RECT 127.075 32.655 127.260 32.745 ;
        RECT 127.850 32.655 128.685 32.665 ;
        RECT 127.075 32.455 128.685 32.655 ;
        RECT 127.075 32.415 127.305 32.455 ;
        RECT 126.570 32.075 126.905 32.295 ;
        RECT 127.910 31.905 128.265 32.285 ;
        RECT 128.435 32.075 128.685 32.455 ;
        RECT 128.935 31.905 129.185 32.685 ;
        RECT 129.355 32.075 129.615 32.755 ;
        RECT 129.785 31.905 130.995 32.995 ;
        RECT 131.165 31.905 131.485 33.085 ;
        RECT 131.655 32.925 131.985 33.095 ;
        RECT 133.490 33.045 133.765 33.645 ;
        RECT 131.655 32.135 131.855 32.925 ;
        RECT 132.155 32.835 133.765 33.045 ;
        RECT 132.155 32.735 132.565 32.835 ;
        RECT 132.180 32.075 132.565 32.735 ;
        RECT 132.960 31.905 133.745 32.665 ;
        RECT 133.935 32.075 134.215 34.175 ;
        RECT 134.385 33.910 139.730 34.455 ;
        RECT 135.970 33.080 136.310 33.910 ;
        RECT 139.905 33.685 142.495 34.455 ;
        RECT 142.665 33.730 142.955 34.455 ;
        RECT 143.125 33.685 145.715 34.455 ;
        RECT 137.790 32.340 138.140 33.590 ;
        RECT 139.905 33.165 141.115 33.685 ;
        RECT 141.285 32.995 142.495 33.515 ;
        RECT 143.125 33.165 144.335 33.685 ;
        RECT 146.365 33.645 146.605 34.455 ;
        RECT 146.775 33.645 147.105 34.285 ;
        RECT 147.275 33.645 147.545 34.455 ;
        RECT 134.385 31.905 139.730 32.340 ;
        RECT 139.905 31.905 142.495 32.995 ;
        RECT 142.665 31.905 142.955 33.070 ;
        RECT 144.505 32.995 145.715 33.515 ;
        RECT 146.345 33.215 146.695 33.465 ;
        RECT 146.865 33.045 147.035 33.645 ;
        RECT 147.765 33.635 147.995 34.455 ;
        RECT 148.165 33.655 148.495 34.285 ;
        RECT 147.205 33.215 147.555 33.465 ;
        RECT 147.745 33.215 148.075 33.465 ;
        RECT 148.245 33.055 148.495 33.655 ;
        RECT 148.665 33.635 148.875 34.455 ;
        RECT 149.565 33.780 149.825 34.285 ;
        RECT 150.005 34.075 150.335 34.455 ;
        RECT 150.515 33.905 150.685 34.285 ;
        RECT 143.125 31.905 145.715 32.995 ;
        RECT 146.355 32.875 147.035 33.045 ;
        RECT 146.355 32.090 146.685 32.875 ;
        RECT 147.215 31.905 147.545 33.045 ;
        RECT 147.765 31.905 147.995 33.045 ;
        RECT 148.165 32.075 148.495 33.055 ;
        RECT 148.665 31.905 148.875 33.045 ;
        RECT 149.565 32.980 149.745 33.780 ;
        RECT 150.020 33.735 150.685 33.905 ;
        RECT 150.020 33.480 150.190 33.735 ;
        RECT 150.945 33.705 152.155 34.455 ;
        RECT 149.915 33.150 150.190 33.480 ;
        RECT 150.415 33.185 150.755 33.555 ;
        RECT 150.020 33.005 150.190 33.150 ;
        RECT 149.565 32.075 149.835 32.980 ;
        RECT 150.020 32.835 150.695 33.005 ;
        RECT 150.005 31.905 150.335 32.665 ;
        RECT 150.515 32.075 150.695 32.835 ;
        RECT 150.945 32.995 151.465 33.535 ;
        RECT 151.635 33.165 152.155 33.705 ;
        RECT 150.945 31.905 152.155 32.995 ;
        RECT 91.060 31.735 152.240 31.905 ;
        RECT 6.030 29.555 6.380 30.940 ;
        RECT 91.145 30.645 92.355 31.735 ;
        RECT 91.145 29.935 91.665 30.475 ;
        RECT 91.835 30.105 92.355 30.645 ;
        RECT 92.605 30.805 92.785 31.565 ;
        RECT 92.965 30.975 93.295 31.735 ;
        RECT 92.605 30.635 93.280 30.805 ;
        RECT 93.465 30.660 93.735 31.565 ;
        RECT 93.110 30.490 93.280 30.635 ;
        RECT 92.545 30.085 92.885 30.455 ;
        RECT 93.110 30.160 93.385 30.490 ;
        RECT 7.855 29.555 8.595 29.690 ;
        RECT 6.025 28.770 8.595 29.555 ;
        RECT 91.145 29.185 92.355 29.935 ;
        RECT 93.110 29.905 93.280 30.160 ;
        RECT 92.615 29.735 93.280 29.905 ;
        RECT 93.555 29.860 93.735 30.660 ;
        RECT 93.905 30.645 97.415 31.735 ;
        RECT 92.615 29.355 92.785 29.735 ;
        RECT 92.965 29.185 93.295 29.565 ;
        RECT 93.475 29.355 93.735 29.860 ;
        RECT 93.905 29.955 95.555 30.475 ;
        RECT 95.725 30.125 97.415 30.645 ;
        RECT 98.585 30.805 98.765 31.565 ;
        RECT 98.945 30.975 99.275 31.735 ;
        RECT 98.585 30.635 99.260 30.805 ;
        RECT 99.445 30.660 99.715 31.565 ;
        RECT 99.090 30.490 99.260 30.635 ;
        RECT 98.525 30.085 98.865 30.455 ;
        RECT 99.090 30.160 99.365 30.490 ;
        RECT 93.905 29.185 97.415 29.955 ;
        RECT 99.090 29.905 99.260 30.160 ;
        RECT 98.595 29.735 99.260 29.905 ;
        RECT 99.535 29.860 99.715 30.660 ;
        RECT 99.885 30.645 103.395 31.735 ;
        RECT 98.595 29.355 98.765 29.735 ;
        RECT 98.945 29.185 99.275 29.565 ;
        RECT 99.455 29.355 99.715 29.860 ;
        RECT 99.885 29.955 101.535 30.475 ;
        RECT 101.705 30.125 103.395 30.645 ;
        RECT 104.025 30.570 104.315 31.735 ;
        RECT 104.485 30.645 106.155 31.735 ;
        RECT 104.485 29.955 105.235 30.475 ;
        RECT 105.405 30.125 106.155 30.645 ;
        RECT 106.405 30.805 106.585 31.565 ;
        RECT 106.765 30.975 107.095 31.735 ;
        RECT 106.405 30.635 107.080 30.805 ;
        RECT 107.265 30.660 107.535 31.565 ;
        RECT 107.705 31.300 113.050 31.735 ;
        RECT 106.910 30.490 107.080 30.635 ;
        RECT 106.345 30.085 106.685 30.455 ;
        RECT 106.910 30.160 107.185 30.490 ;
        RECT 99.885 29.185 103.395 29.955 ;
        RECT 104.025 29.185 104.315 29.910 ;
        RECT 104.485 29.185 106.155 29.955 ;
        RECT 106.910 29.905 107.080 30.160 ;
        RECT 106.415 29.735 107.080 29.905 ;
        RECT 107.355 29.860 107.535 30.660 ;
        RECT 106.415 29.355 106.585 29.735 ;
        RECT 106.765 29.185 107.095 29.565 ;
        RECT 107.275 29.355 107.535 29.860 ;
        RECT 109.290 29.730 109.630 30.560 ;
        RECT 111.110 30.050 111.460 31.300 ;
        RECT 114.225 30.805 114.405 31.565 ;
        RECT 114.585 30.975 114.915 31.735 ;
        RECT 114.225 30.635 114.900 30.805 ;
        RECT 115.085 30.660 115.355 31.565 ;
        RECT 114.730 30.490 114.900 30.635 ;
        RECT 114.165 30.085 114.505 30.455 ;
        RECT 114.730 30.160 115.005 30.490 ;
        RECT 114.730 29.905 114.900 30.160 ;
        RECT 114.235 29.735 114.900 29.905 ;
        RECT 115.175 29.860 115.355 30.660 ;
        RECT 115.525 30.645 116.735 31.735 ;
        RECT 107.705 29.185 113.050 29.730 ;
        RECT 114.235 29.355 114.405 29.735 ;
        RECT 114.585 29.185 114.915 29.565 ;
        RECT 115.095 29.355 115.355 29.860 ;
        RECT 115.525 29.935 116.045 30.475 ;
        RECT 116.215 30.105 116.735 30.645 ;
        RECT 116.905 30.570 117.195 31.735 ;
        RECT 117.365 30.645 118.575 31.735 ;
        RECT 117.365 29.935 117.885 30.475 ;
        RECT 118.055 30.105 118.575 30.645 ;
        RECT 118.805 30.595 119.015 31.735 ;
        RECT 119.185 30.585 119.515 31.565 ;
        RECT 119.685 30.595 119.915 31.735 ;
        RECT 120.125 30.645 121.795 31.735 ;
        RECT 115.525 29.185 116.735 29.935 ;
        RECT 116.905 29.185 117.195 29.910 ;
        RECT 117.365 29.185 118.575 29.935 ;
        RECT 118.805 29.185 119.015 30.005 ;
        RECT 119.185 29.985 119.435 30.585 ;
        RECT 119.605 30.175 119.935 30.425 ;
        RECT 119.185 29.355 119.515 29.985 ;
        RECT 119.685 29.185 119.915 30.005 ;
        RECT 120.125 29.955 120.875 30.475 ;
        RECT 121.045 30.125 121.795 30.645 ;
        RECT 121.965 30.660 122.235 31.565 ;
        RECT 122.405 30.975 122.735 31.735 ;
        RECT 122.915 30.805 123.095 31.565 ;
        RECT 123.345 31.300 128.690 31.735 ;
        RECT 120.125 29.185 121.795 29.955 ;
        RECT 121.965 29.860 122.145 30.660 ;
        RECT 122.420 30.635 123.095 30.805 ;
        RECT 122.420 30.490 122.590 30.635 ;
        RECT 122.315 30.160 122.590 30.490 ;
        RECT 122.420 29.905 122.590 30.160 ;
        RECT 122.815 30.085 123.155 30.455 ;
        RECT 121.965 29.355 122.225 29.860 ;
        RECT 122.420 29.735 123.085 29.905 ;
        RECT 122.405 29.185 122.735 29.565 ;
        RECT 122.915 29.355 123.085 29.735 ;
        RECT 124.930 29.730 125.270 30.560 ;
        RECT 126.750 30.050 127.100 31.300 ;
        RECT 129.785 30.570 130.075 31.735 ;
        RECT 130.245 30.660 130.515 31.565 ;
        RECT 130.685 30.975 131.015 31.735 ;
        RECT 131.195 30.805 131.375 31.565 ;
        RECT 131.625 31.300 136.970 31.735 ;
        RECT 123.345 29.185 128.690 29.730 ;
        RECT 129.785 29.185 130.075 29.910 ;
        RECT 130.245 29.860 130.425 30.660 ;
        RECT 130.700 30.635 131.375 30.805 ;
        RECT 130.700 30.490 130.870 30.635 ;
        RECT 130.595 30.160 130.870 30.490 ;
        RECT 130.700 29.905 130.870 30.160 ;
        RECT 131.095 30.085 131.435 30.455 ;
        RECT 130.245 29.355 130.505 29.860 ;
        RECT 130.700 29.735 131.365 29.905 ;
        RECT 130.685 29.185 131.015 29.565 ;
        RECT 131.195 29.355 131.365 29.735 ;
        RECT 133.210 29.730 133.550 30.560 ;
        RECT 135.030 30.050 135.380 31.300 ;
        RECT 137.605 30.660 137.875 31.565 ;
        RECT 138.045 30.975 138.375 31.735 ;
        RECT 138.555 30.805 138.735 31.565 ;
        RECT 137.605 29.860 137.785 30.660 ;
        RECT 138.060 30.635 138.735 30.805 ;
        RECT 138.985 30.645 142.495 31.735 ;
        RECT 138.060 30.490 138.230 30.635 ;
        RECT 137.955 30.160 138.230 30.490 ;
        RECT 138.060 29.905 138.230 30.160 ;
        RECT 138.455 30.085 138.795 30.455 ;
        RECT 138.985 29.955 140.635 30.475 ;
        RECT 140.805 30.125 142.495 30.645 ;
        RECT 142.665 30.570 142.955 31.735 ;
        RECT 143.125 31.140 143.560 31.565 ;
        RECT 143.730 31.310 144.115 31.735 ;
        RECT 143.125 30.970 144.115 31.140 ;
        RECT 143.125 30.095 143.610 30.800 ;
        RECT 143.780 30.425 144.115 30.970 ;
        RECT 144.285 30.775 144.710 31.565 ;
        RECT 144.880 31.140 145.155 31.565 ;
        RECT 145.325 31.310 145.710 31.735 ;
        RECT 144.880 30.945 145.710 31.140 ;
        RECT 144.285 30.595 145.190 30.775 ;
        RECT 143.780 30.095 144.190 30.425 ;
        RECT 144.360 30.095 145.190 30.595 ;
        RECT 145.360 30.425 145.710 30.945 ;
        RECT 145.880 30.775 146.125 31.565 ;
        RECT 146.315 31.140 146.570 31.565 ;
        RECT 146.740 31.310 147.125 31.735 ;
        RECT 146.315 30.945 147.125 31.140 ;
        RECT 145.880 30.595 146.605 30.775 ;
        RECT 145.360 30.095 145.785 30.425 ;
        RECT 145.955 30.095 146.605 30.595 ;
        RECT 146.775 30.425 147.125 30.945 ;
        RECT 147.295 30.595 147.555 31.565 ;
        RECT 147.725 30.645 148.935 31.735 ;
        RECT 149.110 31.310 149.445 31.735 ;
        RECT 149.615 31.130 149.800 31.535 ;
        RECT 146.775 30.095 147.200 30.425 ;
        RECT 131.625 29.185 136.970 29.730 ;
        RECT 137.605 29.355 137.865 29.860 ;
        RECT 138.060 29.735 138.725 29.905 ;
        RECT 138.045 29.185 138.375 29.565 ;
        RECT 138.555 29.355 138.725 29.735 ;
        RECT 138.985 29.185 142.495 29.955 ;
        RECT 143.780 29.925 144.115 30.095 ;
        RECT 144.360 29.925 144.710 30.095 ;
        RECT 145.360 29.925 145.710 30.095 ;
        RECT 145.955 29.925 146.125 30.095 ;
        RECT 146.775 29.925 147.125 30.095 ;
        RECT 147.370 29.925 147.555 30.595 ;
        RECT 142.665 29.185 142.955 29.910 ;
        RECT 143.125 29.755 144.115 29.925 ;
        RECT 143.125 29.355 143.560 29.755 ;
        RECT 143.730 29.185 144.115 29.585 ;
        RECT 144.285 29.355 144.710 29.925 ;
        RECT 144.900 29.755 145.710 29.925 ;
        RECT 144.900 29.355 145.155 29.755 ;
        RECT 145.325 29.185 145.710 29.585 ;
        RECT 145.880 29.355 146.125 29.925 ;
        RECT 146.315 29.755 147.125 29.925 ;
        RECT 146.315 29.355 146.570 29.755 ;
        RECT 146.740 29.185 147.125 29.585 ;
        RECT 147.295 29.355 147.555 29.925 ;
        RECT 147.725 29.935 148.245 30.475 ;
        RECT 148.415 30.105 148.935 30.645 ;
        RECT 149.135 30.955 149.800 31.130 ;
        RECT 150.005 30.955 150.335 31.735 ;
        RECT 147.725 29.185 148.935 29.935 ;
        RECT 149.135 29.925 149.475 30.955 ;
        RECT 150.505 30.765 150.775 31.535 ;
        RECT 149.645 30.595 150.775 30.765 ;
        RECT 149.645 30.095 149.895 30.595 ;
        RECT 149.135 29.755 149.820 29.925 ;
        RECT 150.075 29.845 150.435 30.425 ;
        RECT 149.110 29.185 149.445 29.585 ;
        RECT 149.615 29.355 149.820 29.755 ;
        RECT 150.605 29.685 150.775 30.595 ;
        RECT 150.945 30.645 152.155 31.735 ;
        RECT 150.945 30.105 151.465 30.645 ;
        RECT 151.635 29.935 152.155 30.475 ;
        RECT 150.030 29.185 150.305 29.665 ;
        RECT 150.515 29.355 150.775 29.685 ;
        RECT 150.945 29.185 152.155 29.935 ;
        RECT 91.060 29.015 152.240 29.185 ;
        RECT 6.030 21.940 6.370 28.770 ;
        RECT 7.855 28.675 8.595 28.770 ;
        RECT 59.055 24.665 59.405 26.505 ;
        RECT 6.020 19.780 6.370 21.940 ;
        RECT 59.050 20.940 59.420 24.665 ;
        RECT 59.010 20.540 59.440 20.940 ;
        RECT 6.020 18.125 6.370 18.780 ;
        RECT 8.230 18.125 10.045 18.735 ;
        RECT 6.020 16.630 10.045 18.125 ;
        RECT 6.020 16.620 6.370 16.630 ;
        RECT 8.230 15.990 10.045 16.630 ;
        RECT 59.050 12.320 59.420 20.540 ;
        RECT 59.060 10.430 59.410 12.320 ;
        RECT 59.060 8.675 59.410 9.930 ;
        RECT 53.125 7.780 59.410 8.675 ;
        RECT 59.060 7.770 59.410 7.780 ;
      LAYER mcon ;
        RECT 71.395 194.345 71.565 194.515 ;
        RECT 71.855 194.345 72.025 194.515 ;
        RECT 72.315 194.345 72.485 194.515 ;
        RECT 72.775 194.345 72.945 194.515 ;
        RECT 73.235 194.345 73.405 194.515 ;
        RECT 73.695 194.345 73.865 194.515 ;
        RECT 74.155 194.345 74.325 194.515 ;
        RECT 74.615 194.345 74.785 194.515 ;
        RECT 75.075 194.345 75.245 194.515 ;
        RECT 75.535 194.345 75.705 194.515 ;
        RECT 75.995 194.345 76.165 194.515 ;
        RECT 76.455 194.345 76.625 194.515 ;
        RECT 76.915 194.345 77.085 194.515 ;
        RECT 77.375 194.345 77.545 194.515 ;
        RECT 77.835 194.345 78.005 194.515 ;
        RECT 78.295 194.345 78.465 194.515 ;
        RECT 78.755 194.345 78.925 194.515 ;
        RECT 79.215 194.345 79.385 194.515 ;
        RECT 79.675 194.345 79.845 194.515 ;
        RECT 80.135 194.345 80.305 194.515 ;
        RECT 80.595 194.345 80.765 194.515 ;
        RECT 81.055 194.345 81.225 194.515 ;
        RECT 81.515 194.345 81.685 194.515 ;
        RECT 81.975 194.345 82.145 194.515 ;
        RECT 82.435 194.345 82.605 194.515 ;
        RECT 82.895 194.345 83.065 194.515 ;
        RECT 83.355 194.345 83.525 194.515 ;
        RECT 83.815 194.345 83.985 194.515 ;
        RECT 84.275 194.345 84.445 194.515 ;
        RECT 84.735 194.345 84.905 194.515 ;
        RECT 85.195 194.345 85.365 194.515 ;
        RECT 85.655 194.345 85.825 194.515 ;
        RECT 86.115 194.345 86.285 194.515 ;
        RECT 86.575 194.345 86.745 194.515 ;
        RECT 87.035 194.345 87.205 194.515 ;
        RECT 87.495 194.345 87.665 194.515 ;
        RECT 87.955 194.345 88.125 194.515 ;
        RECT 88.415 194.345 88.585 194.515 ;
        RECT 88.875 194.345 89.045 194.515 ;
        RECT 89.335 194.345 89.505 194.515 ;
        RECT 89.795 194.345 89.965 194.515 ;
        RECT 90.255 194.345 90.425 194.515 ;
        RECT 90.715 194.345 90.885 194.515 ;
        RECT 91.175 194.345 91.345 194.515 ;
        RECT 91.635 194.345 91.805 194.515 ;
        RECT 92.095 194.345 92.265 194.515 ;
        RECT 92.555 194.345 92.725 194.515 ;
        RECT 93.015 194.345 93.185 194.515 ;
        RECT 93.475 194.345 93.645 194.515 ;
        RECT 93.935 194.345 94.105 194.515 ;
        RECT 94.395 194.345 94.565 194.515 ;
        RECT 94.855 194.345 95.025 194.515 ;
        RECT 95.315 194.345 95.485 194.515 ;
        RECT 95.775 194.345 95.945 194.515 ;
        RECT 96.235 194.345 96.405 194.515 ;
        RECT 96.695 194.345 96.865 194.515 ;
        RECT 97.155 194.345 97.325 194.515 ;
        RECT 97.615 194.345 97.785 194.515 ;
        RECT 98.075 194.345 98.245 194.515 ;
        RECT 98.535 194.345 98.705 194.515 ;
        RECT 98.995 194.345 99.165 194.515 ;
        RECT 99.455 194.345 99.625 194.515 ;
        RECT 99.915 194.345 100.085 194.515 ;
        RECT 100.375 194.345 100.545 194.515 ;
        RECT 100.835 194.345 101.005 194.515 ;
        RECT 101.295 194.345 101.465 194.515 ;
        RECT 101.755 194.345 101.925 194.515 ;
        RECT 102.215 194.345 102.385 194.515 ;
        RECT 102.675 194.345 102.845 194.515 ;
        RECT 103.135 194.345 103.305 194.515 ;
        RECT 103.595 194.345 103.765 194.515 ;
        RECT 104.055 194.345 104.225 194.515 ;
        RECT 104.515 194.345 104.685 194.515 ;
        RECT 104.975 194.345 105.145 194.515 ;
        RECT 105.435 194.345 105.605 194.515 ;
        RECT 105.895 194.345 106.065 194.515 ;
        RECT 106.355 194.345 106.525 194.515 ;
        RECT 106.815 194.345 106.985 194.515 ;
        RECT 107.275 194.345 107.445 194.515 ;
        RECT 107.735 194.345 107.905 194.515 ;
        RECT 108.195 194.345 108.365 194.515 ;
        RECT 108.655 194.345 108.825 194.515 ;
        RECT 109.115 194.345 109.285 194.515 ;
        RECT 109.575 194.345 109.745 194.515 ;
        RECT 110.035 194.345 110.205 194.515 ;
        RECT 110.495 194.345 110.665 194.515 ;
        RECT 110.955 194.345 111.125 194.515 ;
        RECT 111.415 194.345 111.585 194.515 ;
        RECT 111.875 194.345 112.045 194.515 ;
        RECT 112.335 194.345 112.505 194.515 ;
        RECT 112.795 194.345 112.965 194.515 ;
        RECT 113.255 194.345 113.425 194.515 ;
        RECT 113.715 194.345 113.885 194.515 ;
        RECT 114.175 194.345 114.345 194.515 ;
        RECT 114.635 194.345 114.805 194.515 ;
        RECT 115.095 194.345 115.265 194.515 ;
        RECT 115.555 194.345 115.725 194.515 ;
        RECT 116.015 194.345 116.185 194.515 ;
        RECT 116.475 194.345 116.645 194.515 ;
        RECT 116.935 194.345 117.105 194.515 ;
        RECT 117.395 194.345 117.565 194.515 ;
        RECT 117.855 194.345 118.025 194.515 ;
        RECT 118.315 194.345 118.485 194.515 ;
        RECT 118.775 194.345 118.945 194.515 ;
        RECT 119.235 194.345 119.405 194.515 ;
        RECT 81.975 193.835 82.145 194.005 ;
        RECT 81.515 192.475 81.685 192.645 ;
        RECT 86.115 192.135 86.285 192.305 ;
        RECT 88.875 192.815 89.045 192.985 ;
        RECT 101.295 192.475 101.465 192.645 ;
        RECT 111.875 193.835 112.045 194.005 ;
        RECT 102.215 192.135 102.385 192.305 ;
        RECT 111.415 192.475 111.585 192.645 ;
        RECT 71.395 191.625 71.565 191.795 ;
        RECT 71.855 191.625 72.025 191.795 ;
        RECT 72.315 191.625 72.485 191.795 ;
        RECT 72.775 191.625 72.945 191.795 ;
        RECT 73.235 191.625 73.405 191.795 ;
        RECT 73.695 191.625 73.865 191.795 ;
        RECT 74.155 191.625 74.325 191.795 ;
        RECT 74.615 191.625 74.785 191.795 ;
        RECT 75.075 191.625 75.245 191.795 ;
        RECT 75.535 191.625 75.705 191.795 ;
        RECT 75.995 191.625 76.165 191.795 ;
        RECT 76.455 191.625 76.625 191.795 ;
        RECT 76.915 191.625 77.085 191.795 ;
        RECT 77.375 191.625 77.545 191.795 ;
        RECT 77.835 191.625 78.005 191.795 ;
        RECT 78.295 191.625 78.465 191.795 ;
        RECT 78.755 191.625 78.925 191.795 ;
        RECT 79.215 191.625 79.385 191.795 ;
        RECT 79.675 191.625 79.845 191.795 ;
        RECT 80.135 191.625 80.305 191.795 ;
        RECT 80.595 191.625 80.765 191.795 ;
        RECT 81.055 191.625 81.225 191.795 ;
        RECT 81.515 191.625 81.685 191.795 ;
        RECT 81.975 191.625 82.145 191.795 ;
        RECT 82.435 191.625 82.605 191.795 ;
        RECT 82.895 191.625 83.065 191.795 ;
        RECT 83.355 191.625 83.525 191.795 ;
        RECT 83.815 191.625 83.985 191.795 ;
        RECT 84.275 191.625 84.445 191.795 ;
        RECT 84.735 191.625 84.905 191.795 ;
        RECT 85.195 191.625 85.365 191.795 ;
        RECT 85.655 191.625 85.825 191.795 ;
        RECT 86.115 191.625 86.285 191.795 ;
        RECT 86.575 191.625 86.745 191.795 ;
        RECT 87.035 191.625 87.205 191.795 ;
        RECT 87.495 191.625 87.665 191.795 ;
        RECT 87.955 191.625 88.125 191.795 ;
        RECT 88.415 191.625 88.585 191.795 ;
        RECT 88.875 191.625 89.045 191.795 ;
        RECT 89.335 191.625 89.505 191.795 ;
        RECT 89.795 191.625 89.965 191.795 ;
        RECT 90.255 191.625 90.425 191.795 ;
        RECT 90.715 191.625 90.885 191.795 ;
        RECT 91.175 191.625 91.345 191.795 ;
        RECT 91.635 191.625 91.805 191.795 ;
        RECT 92.095 191.625 92.265 191.795 ;
        RECT 92.555 191.625 92.725 191.795 ;
        RECT 93.015 191.625 93.185 191.795 ;
        RECT 93.475 191.625 93.645 191.795 ;
        RECT 93.935 191.625 94.105 191.795 ;
        RECT 94.395 191.625 94.565 191.795 ;
        RECT 94.855 191.625 95.025 191.795 ;
        RECT 95.315 191.625 95.485 191.795 ;
        RECT 95.775 191.625 95.945 191.795 ;
        RECT 96.235 191.625 96.405 191.795 ;
        RECT 96.695 191.625 96.865 191.795 ;
        RECT 97.155 191.625 97.325 191.795 ;
        RECT 97.615 191.625 97.785 191.795 ;
        RECT 98.075 191.625 98.245 191.795 ;
        RECT 98.535 191.625 98.705 191.795 ;
        RECT 98.995 191.625 99.165 191.795 ;
        RECT 99.455 191.625 99.625 191.795 ;
        RECT 99.915 191.625 100.085 191.795 ;
        RECT 100.375 191.625 100.545 191.795 ;
        RECT 100.835 191.625 101.005 191.795 ;
        RECT 101.295 191.625 101.465 191.795 ;
        RECT 101.755 191.625 101.925 191.795 ;
        RECT 102.215 191.625 102.385 191.795 ;
        RECT 102.675 191.625 102.845 191.795 ;
        RECT 103.135 191.625 103.305 191.795 ;
        RECT 103.595 191.625 103.765 191.795 ;
        RECT 104.055 191.625 104.225 191.795 ;
        RECT 104.515 191.625 104.685 191.795 ;
        RECT 104.975 191.625 105.145 191.795 ;
        RECT 105.435 191.625 105.605 191.795 ;
        RECT 105.895 191.625 106.065 191.795 ;
        RECT 106.355 191.625 106.525 191.795 ;
        RECT 106.815 191.625 106.985 191.795 ;
        RECT 107.275 191.625 107.445 191.795 ;
        RECT 107.735 191.625 107.905 191.795 ;
        RECT 108.195 191.625 108.365 191.795 ;
        RECT 108.655 191.625 108.825 191.795 ;
        RECT 109.115 191.625 109.285 191.795 ;
        RECT 109.575 191.625 109.745 191.795 ;
        RECT 110.035 191.625 110.205 191.795 ;
        RECT 110.495 191.625 110.665 191.795 ;
        RECT 110.955 191.625 111.125 191.795 ;
        RECT 111.415 191.625 111.585 191.795 ;
        RECT 111.875 191.625 112.045 191.795 ;
        RECT 112.335 191.625 112.505 191.795 ;
        RECT 112.795 191.625 112.965 191.795 ;
        RECT 113.255 191.625 113.425 191.795 ;
        RECT 113.715 191.625 113.885 191.795 ;
        RECT 114.175 191.625 114.345 191.795 ;
        RECT 114.635 191.625 114.805 191.795 ;
        RECT 115.095 191.625 115.265 191.795 ;
        RECT 115.555 191.625 115.725 191.795 ;
        RECT 116.015 191.625 116.185 191.795 ;
        RECT 116.475 191.625 116.645 191.795 ;
        RECT 116.935 191.625 117.105 191.795 ;
        RECT 117.395 191.625 117.565 191.795 ;
        RECT 117.855 191.625 118.025 191.795 ;
        RECT 118.315 191.625 118.485 191.795 ;
        RECT 118.775 191.625 118.945 191.795 ;
        RECT 119.235 191.625 119.405 191.795 ;
        RECT 72.775 190.435 72.945 190.605 ;
        RECT 77.375 191.115 77.545 191.285 ;
        RECT 73.695 189.415 73.865 189.585 ;
        RECT 79.630 190.095 79.800 190.265 ;
        RECT 81.055 190.435 81.225 190.605 ;
        RECT 80.135 189.755 80.305 189.925 ;
        RECT 81.510 189.755 81.680 189.925 ;
        RECT 81.970 190.095 82.140 190.265 ;
        RECT 82.895 190.435 83.065 190.605 ;
        RECT 82.435 190.095 82.605 190.265 ;
        RECT 83.815 190.435 83.985 190.605 ;
        RECT 83.355 189.415 83.525 189.585 ;
        RECT 87.035 189.415 87.205 189.585 ;
        RECT 89.345 190.095 89.515 190.265 ;
        RECT 89.780 189.755 89.950 189.925 ;
        RECT 91.865 190.095 92.035 190.265 ;
        RECT 91.350 189.755 91.520 189.925 ;
        RECT 92.710 190.775 92.880 190.945 ;
        RECT 93.055 190.095 93.225 190.265 ;
        RECT 93.935 190.095 94.105 190.265 ;
        RECT 94.395 190.095 94.565 190.265 ;
        RECT 95.315 190.435 95.485 190.605 ;
        RECT 95.775 190.435 95.945 190.605 ;
        RECT 93.450 189.755 93.620 189.925 ;
        RECT 97.615 189.415 97.785 189.585 ;
        RECT 100.835 190.095 101.005 190.265 ;
        RECT 102.215 190.435 102.385 190.605 ;
        RECT 103.135 190.435 103.305 190.605 ;
        RECT 103.595 190.435 103.765 190.605 ;
        RECT 101.295 189.755 101.465 189.925 ;
        RECT 105.895 190.435 106.065 190.605 ;
        RECT 106.360 190.095 106.530 190.265 ;
        RECT 107.275 190.435 107.445 190.605 ;
        RECT 106.820 189.755 106.990 189.925 ;
        RECT 108.195 189.755 108.365 189.925 ;
        RECT 108.700 190.095 108.870 190.265 ;
        RECT 110.955 191.115 111.125 191.285 ;
        RECT 117.855 190.435 118.025 190.605 ;
        RECT 116.935 189.415 117.105 189.585 ;
        RECT 71.395 188.905 71.565 189.075 ;
        RECT 71.855 188.905 72.025 189.075 ;
        RECT 72.315 188.905 72.485 189.075 ;
        RECT 72.775 188.905 72.945 189.075 ;
        RECT 73.235 188.905 73.405 189.075 ;
        RECT 73.695 188.905 73.865 189.075 ;
        RECT 74.155 188.905 74.325 189.075 ;
        RECT 74.615 188.905 74.785 189.075 ;
        RECT 75.075 188.905 75.245 189.075 ;
        RECT 75.535 188.905 75.705 189.075 ;
        RECT 75.995 188.905 76.165 189.075 ;
        RECT 76.455 188.905 76.625 189.075 ;
        RECT 76.915 188.905 77.085 189.075 ;
        RECT 77.375 188.905 77.545 189.075 ;
        RECT 77.835 188.905 78.005 189.075 ;
        RECT 78.295 188.905 78.465 189.075 ;
        RECT 78.755 188.905 78.925 189.075 ;
        RECT 79.215 188.905 79.385 189.075 ;
        RECT 79.675 188.905 79.845 189.075 ;
        RECT 80.135 188.905 80.305 189.075 ;
        RECT 80.595 188.905 80.765 189.075 ;
        RECT 81.055 188.905 81.225 189.075 ;
        RECT 81.515 188.905 81.685 189.075 ;
        RECT 81.975 188.905 82.145 189.075 ;
        RECT 82.435 188.905 82.605 189.075 ;
        RECT 82.895 188.905 83.065 189.075 ;
        RECT 83.355 188.905 83.525 189.075 ;
        RECT 83.815 188.905 83.985 189.075 ;
        RECT 84.275 188.905 84.445 189.075 ;
        RECT 84.735 188.905 84.905 189.075 ;
        RECT 85.195 188.905 85.365 189.075 ;
        RECT 85.655 188.905 85.825 189.075 ;
        RECT 86.115 188.905 86.285 189.075 ;
        RECT 86.575 188.905 86.745 189.075 ;
        RECT 87.035 188.905 87.205 189.075 ;
        RECT 87.495 188.905 87.665 189.075 ;
        RECT 87.955 188.905 88.125 189.075 ;
        RECT 88.415 188.905 88.585 189.075 ;
        RECT 88.875 188.905 89.045 189.075 ;
        RECT 89.335 188.905 89.505 189.075 ;
        RECT 89.795 188.905 89.965 189.075 ;
        RECT 90.255 188.905 90.425 189.075 ;
        RECT 90.715 188.905 90.885 189.075 ;
        RECT 91.175 188.905 91.345 189.075 ;
        RECT 91.635 188.905 91.805 189.075 ;
        RECT 92.095 188.905 92.265 189.075 ;
        RECT 92.555 188.905 92.725 189.075 ;
        RECT 93.015 188.905 93.185 189.075 ;
        RECT 93.475 188.905 93.645 189.075 ;
        RECT 93.935 188.905 94.105 189.075 ;
        RECT 94.395 188.905 94.565 189.075 ;
        RECT 94.855 188.905 95.025 189.075 ;
        RECT 95.315 188.905 95.485 189.075 ;
        RECT 95.775 188.905 95.945 189.075 ;
        RECT 96.235 188.905 96.405 189.075 ;
        RECT 96.695 188.905 96.865 189.075 ;
        RECT 97.155 188.905 97.325 189.075 ;
        RECT 97.615 188.905 97.785 189.075 ;
        RECT 98.075 188.905 98.245 189.075 ;
        RECT 98.535 188.905 98.705 189.075 ;
        RECT 98.995 188.905 99.165 189.075 ;
        RECT 99.455 188.905 99.625 189.075 ;
        RECT 99.915 188.905 100.085 189.075 ;
        RECT 100.375 188.905 100.545 189.075 ;
        RECT 100.835 188.905 101.005 189.075 ;
        RECT 101.295 188.905 101.465 189.075 ;
        RECT 101.755 188.905 101.925 189.075 ;
        RECT 102.215 188.905 102.385 189.075 ;
        RECT 102.675 188.905 102.845 189.075 ;
        RECT 103.135 188.905 103.305 189.075 ;
        RECT 103.595 188.905 103.765 189.075 ;
        RECT 104.055 188.905 104.225 189.075 ;
        RECT 104.515 188.905 104.685 189.075 ;
        RECT 104.975 188.905 105.145 189.075 ;
        RECT 105.435 188.905 105.605 189.075 ;
        RECT 105.895 188.905 106.065 189.075 ;
        RECT 106.355 188.905 106.525 189.075 ;
        RECT 106.815 188.905 106.985 189.075 ;
        RECT 107.275 188.905 107.445 189.075 ;
        RECT 107.735 188.905 107.905 189.075 ;
        RECT 108.195 188.905 108.365 189.075 ;
        RECT 108.655 188.905 108.825 189.075 ;
        RECT 109.115 188.905 109.285 189.075 ;
        RECT 109.575 188.905 109.745 189.075 ;
        RECT 110.035 188.905 110.205 189.075 ;
        RECT 110.495 188.905 110.665 189.075 ;
        RECT 110.955 188.905 111.125 189.075 ;
        RECT 111.415 188.905 111.585 189.075 ;
        RECT 111.875 188.905 112.045 189.075 ;
        RECT 112.335 188.905 112.505 189.075 ;
        RECT 112.795 188.905 112.965 189.075 ;
        RECT 113.255 188.905 113.425 189.075 ;
        RECT 113.715 188.905 113.885 189.075 ;
        RECT 114.175 188.905 114.345 189.075 ;
        RECT 114.635 188.905 114.805 189.075 ;
        RECT 115.095 188.905 115.265 189.075 ;
        RECT 115.555 188.905 115.725 189.075 ;
        RECT 116.015 188.905 116.185 189.075 ;
        RECT 116.475 188.905 116.645 189.075 ;
        RECT 116.935 188.905 117.105 189.075 ;
        RECT 117.395 188.905 117.565 189.075 ;
        RECT 117.855 188.905 118.025 189.075 ;
        RECT 118.315 188.905 118.485 189.075 ;
        RECT 118.775 188.905 118.945 189.075 ;
        RECT 119.235 188.905 119.405 189.075 ;
        RECT 82.435 188.395 82.605 188.565 ;
        RECT 83.815 188.395 83.985 188.565 ;
        RECT 82.435 187.715 82.605 187.885 ;
        RECT 80.595 187.375 80.765 187.545 ;
        RECT 82.880 187.375 83.050 187.545 ;
        RECT 85.220 188.055 85.390 188.225 ;
        RECT 84.735 187.715 84.905 187.885 ;
        RECT 85.615 187.715 85.785 187.885 ;
        RECT 85.960 187.035 86.130 187.205 ;
        RECT 87.320 188.055 87.490 188.225 ;
        RECT 86.805 187.715 86.975 187.885 ;
        RECT 88.890 188.055 89.060 188.225 ;
        RECT 89.325 187.715 89.495 187.885 ;
        RECT 92.095 187.035 92.265 187.205 ;
        RECT 91.635 186.695 91.805 186.865 ;
        RECT 97.640 188.055 97.810 188.225 ;
        RECT 94.855 187.375 95.025 187.545 ;
        RECT 95.775 187.375 95.945 187.545 ;
        RECT 97.155 187.715 97.325 187.885 ;
        RECT 96.235 186.695 96.405 186.865 ;
        RECT 98.035 187.715 98.205 187.885 ;
        RECT 98.490 187.035 98.660 187.205 ;
        RECT 99.740 188.055 99.910 188.225 ;
        RECT 99.225 187.715 99.395 187.885 ;
        RECT 101.310 188.055 101.480 188.225 ;
        RECT 101.745 187.715 101.915 187.885 ;
        RECT 104.055 188.395 104.225 188.565 ;
        RECT 105.895 187.715 106.065 187.885 ;
        RECT 105.435 187.375 105.605 187.545 ;
        RECT 106.355 188.055 106.525 188.225 ;
        RECT 107.735 188.395 107.905 188.565 ;
        RECT 106.815 187.375 106.985 187.545 ;
        RECT 104.515 187.035 104.685 187.205 ;
        RECT 107.735 187.375 107.905 187.545 ;
        RECT 112.795 188.395 112.965 188.565 ;
        RECT 108.655 187.375 108.825 187.545 ;
        RECT 111.415 187.375 111.585 187.545 ;
        RECT 115.095 187.375 115.265 187.545 ;
        RECT 114.175 186.695 114.345 186.865 ;
        RECT 71.395 186.185 71.565 186.355 ;
        RECT 71.855 186.185 72.025 186.355 ;
        RECT 72.315 186.185 72.485 186.355 ;
        RECT 72.775 186.185 72.945 186.355 ;
        RECT 73.235 186.185 73.405 186.355 ;
        RECT 73.695 186.185 73.865 186.355 ;
        RECT 74.155 186.185 74.325 186.355 ;
        RECT 74.615 186.185 74.785 186.355 ;
        RECT 75.075 186.185 75.245 186.355 ;
        RECT 75.535 186.185 75.705 186.355 ;
        RECT 75.995 186.185 76.165 186.355 ;
        RECT 76.455 186.185 76.625 186.355 ;
        RECT 76.915 186.185 77.085 186.355 ;
        RECT 77.375 186.185 77.545 186.355 ;
        RECT 77.835 186.185 78.005 186.355 ;
        RECT 78.295 186.185 78.465 186.355 ;
        RECT 78.755 186.185 78.925 186.355 ;
        RECT 79.215 186.185 79.385 186.355 ;
        RECT 79.675 186.185 79.845 186.355 ;
        RECT 80.135 186.185 80.305 186.355 ;
        RECT 80.595 186.185 80.765 186.355 ;
        RECT 81.055 186.185 81.225 186.355 ;
        RECT 81.515 186.185 81.685 186.355 ;
        RECT 81.975 186.185 82.145 186.355 ;
        RECT 82.435 186.185 82.605 186.355 ;
        RECT 82.895 186.185 83.065 186.355 ;
        RECT 83.355 186.185 83.525 186.355 ;
        RECT 83.815 186.185 83.985 186.355 ;
        RECT 84.275 186.185 84.445 186.355 ;
        RECT 84.735 186.185 84.905 186.355 ;
        RECT 85.195 186.185 85.365 186.355 ;
        RECT 85.655 186.185 85.825 186.355 ;
        RECT 86.115 186.185 86.285 186.355 ;
        RECT 86.575 186.185 86.745 186.355 ;
        RECT 87.035 186.185 87.205 186.355 ;
        RECT 87.495 186.185 87.665 186.355 ;
        RECT 87.955 186.185 88.125 186.355 ;
        RECT 88.415 186.185 88.585 186.355 ;
        RECT 88.875 186.185 89.045 186.355 ;
        RECT 89.335 186.185 89.505 186.355 ;
        RECT 89.795 186.185 89.965 186.355 ;
        RECT 90.255 186.185 90.425 186.355 ;
        RECT 90.715 186.185 90.885 186.355 ;
        RECT 91.175 186.185 91.345 186.355 ;
        RECT 91.635 186.185 91.805 186.355 ;
        RECT 92.095 186.185 92.265 186.355 ;
        RECT 92.555 186.185 92.725 186.355 ;
        RECT 93.015 186.185 93.185 186.355 ;
        RECT 93.475 186.185 93.645 186.355 ;
        RECT 93.935 186.185 94.105 186.355 ;
        RECT 94.395 186.185 94.565 186.355 ;
        RECT 94.855 186.185 95.025 186.355 ;
        RECT 95.315 186.185 95.485 186.355 ;
        RECT 95.775 186.185 95.945 186.355 ;
        RECT 96.235 186.185 96.405 186.355 ;
        RECT 96.695 186.185 96.865 186.355 ;
        RECT 97.155 186.185 97.325 186.355 ;
        RECT 97.615 186.185 97.785 186.355 ;
        RECT 98.075 186.185 98.245 186.355 ;
        RECT 98.535 186.185 98.705 186.355 ;
        RECT 98.995 186.185 99.165 186.355 ;
        RECT 99.455 186.185 99.625 186.355 ;
        RECT 99.915 186.185 100.085 186.355 ;
        RECT 100.375 186.185 100.545 186.355 ;
        RECT 100.835 186.185 101.005 186.355 ;
        RECT 101.295 186.185 101.465 186.355 ;
        RECT 101.755 186.185 101.925 186.355 ;
        RECT 102.215 186.185 102.385 186.355 ;
        RECT 102.675 186.185 102.845 186.355 ;
        RECT 103.135 186.185 103.305 186.355 ;
        RECT 103.595 186.185 103.765 186.355 ;
        RECT 104.055 186.185 104.225 186.355 ;
        RECT 104.515 186.185 104.685 186.355 ;
        RECT 104.975 186.185 105.145 186.355 ;
        RECT 105.435 186.185 105.605 186.355 ;
        RECT 105.895 186.185 106.065 186.355 ;
        RECT 106.355 186.185 106.525 186.355 ;
        RECT 106.815 186.185 106.985 186.355 ;
        RECT 107.275 186.185 107.445 186.355 ;
        RECT 107.735 186.185 107.905 186.355 ;
        RECT 108.195 186.185 108.365 186.355 ;
        RECT 108.655 186.185 108.825 186.355 ;
        RECT 109.115 186.185 109.285 186.355 ;
        RECT 109.575 186.185 109.745 186.355 ;
        RECT 110.035 186.185 110.205 186.355 ;
        RECT 110.495 186.185 110.665 186.355 ;
        RECT 110.955 186.185 111.125 186.355 ;
        RECT 111.415 186.185 111.585 186.355 ;
        RECT 111.875 186.185 112.045 186.355 ;
        RECT 112.335 186.185 112.505 186.355 ;
        RECT 112.795 186.185 112.965 186.355 ;
        RECT 113.255 186.185 113.425 186.355 ;
        RECT 113.715 186.185 113.885 186.355 ;
        RECT 114.175 186.185 114.345 186.355 ;
        RECT 114.635 186.185 114.805 186.355 ;
        RECT 115.095 186.185 115.265 186.355 ;
        RECT 115.555 186.185 115.725 186.355 ;
        RECT 116.015 186.185 116.185 186.355 ;
        RECT 116.475 186.185 116.645 186.355 ;
        RECT 116.935 186.185 117.105 186.355 ;
        RECT 117.395 186.185 117.565 186.355 ;
        RECT 117.855 186.185 118.025 186.355 ;
        RECT 118.315 186.185 118.485 186.355 ;
        RECT 118.775 186.185 118.945 186.355 ;
        RECT 119.235 186.185 119.405 186.355 ;
        RECT 85.195 184.995 85.365 185.165 ;
        RECT 86.575 184.995 86.745 185.165 ;
        RECT 83.815 183.975 83.985 184.145 ;
        RECT 86.115 183.975 86.285 184.145 ;
        RECT 89.795 184.655 89.965 184.825 ;
        RECT 91.175 184.655 91.345 184.825 ;
        RECT 93.935 184.655 94.105 184.825 ;
        RECT 98.535 185.675 98.705 185.845 ;
        RECT 96.695 183.975 96.865 184.145 ;
        RECT 99.440 184.995 99.610 185.165 ;
        RECT 104.055 185.675 104.225 185.845 ;
        RECT 102.215 184.995 102.385 185.165 ;
        RECT 102.675 184.995 102.845 185.165 ;
        RECT 101.755 184.655 101.925 184.825 ;
        RECT 101.295 184.315 101.465 184.485 ;
        RECT 102.215 183.975 102.385 184.145 ;
        RECT 107.275 184.995 107.445 185.165 ;
        RECT 106.355 183.975 106.525 184.145 ;
        RECT 108.655 184.995 108.825 185.165 ;
        RECT 107.735 184.315 107.905 184.485 ;
        RECT 110.955 184.655 111.125 184.825 ;
        RECT 111.440 184.315 111.610 184.485 ;
        RECT 111.835 184.655 112.005 184.825 ;
        RECT 112.290 185.335 112.460 185.505 ;
        RECT 113.025 184.655 113.195 184.825 ;
        RECT 113.540 184.315 113.710 184.485 ;
        RECT 115.110 184.315 115.280 184.485 ;
        RECT 115.545 184.655 115.715 184.825 ;
        RECT 117.855 183.975 118.025 184.145 ;
        RECT 71.395 183.465 71.565 183.635 ;
        RECT 71.855 183.465 72.025 183.635 ;
        RECT 72.315 183.465 72.485 183.635 ;
        RECT 72.775 183.465 72.945 183.635 ;
        RECT 73.235 183.465 73.405 183.635 ;
        RECT 73.695 183.465 73.865 183.635 ;
        RECT 74.155 183.465 74.325 183.635 ;
        RECT 74.615 183.465 74.785 183.635 ;
        RECT 75.075 183.465 75.245 183.635 ;
        RECT 75.535 183.465 75.705 183.635 ;
        RECT 75.995 183.465 76.165 183.635 ;
        RECT 76.455 183.465 76.625 183.635 ;
        RECT 76.915 183.465 77.085 183.635 ;
        RECT 77.375 183.465 77.545 183.635 ;
        RECT 77.835 183.465 78.005 183.635 ;
        RECT 78.295 183.465 78.465 183.635 ;
        RECT 78.755 183.465 78.925 183.635 ;
        RECT 79.215 183.465 79.385 183.635 ;
        RECT 79.675 183.465 79.845 183.635 ;
        RECT 80.135 183.465 80.305 183.635 ;
        RECT 80.595 183.465 80.765 183.635 ;
        RECT 81.055 183.465 81.225 183.635 ;
        RECT 81.515 183.465 81.685 183.635 ;
        RECT 81.975 183.465 82.145 183.635 ;
        RECT 82.435 183.465 82.605 183.635 ;
        RECT 82.895 183.465 83.065 183.635 ;
        RECT 83.355 183.465 83.525 183.635 ;
        RECT 83.815 183.465 83.985 183.635 ;
        RECT 84.275 183.465 84.445 183.635 ;
        RECT 84.735 183.465 84.905 183.635 ;
        RECT 85.195 183.465 85.365 183.635 ;
        RECT 85.655 183.465 85.825 183.635 ;
        RECT 86.115 183.465 86.285 183.635 ;
        RECT 86.575 183.465 86.745 183.635 ;
        RECT 87.035 183.465 87.205 183.635 ;
        RECT 87.495 183.465 87.665 183.635 ;
        RECT 87.955 183.465 88.125 183.635 ;
        RECT 88.415 183.465 88.585 183.635 ;
        RECT 88.875 183.465 89.045 183.635 ;
        RECT 89.335 183.465 89.505 183.635 ;
        RECT 89.795 183.465 89.965 183.635 ;
        RECT 90.255 183.465 90.425 183.635 ;
        RECT 90.715 183.465 90.885 183.635 ;
        RECT 91.175 183.465 91.345 183.635 ;
        RECT 91.635 183.465 91.805 183.635 ;
        RECT 92.095 183.465 92.265 183.635 ;
        RECT 92.555 183.465 92.725 183.635 ;
        RECT 93.015 183.465 93.185 183.635 ;
        RECT 93.475 183.465 93.645 183.635 ;
        RECT 93.935 183.465 94.105 183.635 ;
        RECT 94.395 183.465 94.565 183.635 ;
        RECT 94.855 183.465 95.025 183.635 ;
        RECT 95.315 183.465 95.485 183.635 ;
        RECT 95.775 183.465 95.945 183.635 ;
        RECT 96.235 183.465 96.405 183.635 ;
        RECT 96.695 183.465 96.865 183.635 ;
        RECT 97.155 183.465 97.325 183.635 ;
        RECT 97.615 183.465 97.785 183.635 ;
        RECT 98.075 183.465 98.245 183.635 ;
        RECT 98.535 183.465 98.705 183.635 ;
        RECT 98.995 183.465 99.165 183.635 ;
        RECT 99.455 183.465 99.625 183.635 ;
        RECT 99.915 183.465 100.085 183.635 ;
        RECT 100.375 183.465 100.545 183.635 ;
        RECT 100.835 183.465 101.005 183.635 ;
        RECT 101.295 183.465 101.465 183.635 ;
        RECT 101.755 183.465 101.925 183.635 ;
        RECT 102.215 183.465 102.385 183.635 ;
        RECT 102.675 183.465 102.845 183.635 ;
        RECT 103.135 183.465 103.305 183.635 ;
        RECT 103.595 183.465 103.765 183.635 ;
        RECT 104.055 183.465 104.225 183.635 ;
        RECT 104.515 183.465 104.685 183.635 ;
        RECT 104.975 183.465 105.145 183.635 ;
        RECT 105.435 183.465 105.605 183.635 ;
        RECT 105.895 183.465 106.065 183.635 ;
        RECT 106.355 183.465 106.525 183.635 ;
        RECT 106.815 183.465 106.985 183.635 ;
        RECT 107.275 183.465 107.445 183.635 ;
        RECT 107.735 183.465 107.905 183.635 ;
        RECT 108.195 183.465 108.365 183.635 ;
        RECT 108.655 183.465 108.825 183.635 ;
        RECT 109.115 183.465 109.285 183.635 ;
        RECT 109.575 183.465 109.745 183.635 ;
        RECT 110.035 183.465 110.205 183.635 ;
        RECT 110.495 183.465 110.665 183.635 ;
        RECT 110.955 183.465 111.125 183.635 ;
        RECT 111.415 183.465 111.585 183.635 ;
        RECT 111.875 183.465 112.045 183.635 ;
        RECT 112.335 183.465 112.505 183.635 ;
        RECT 112.795 183.465 112.965 183.635 ;
        RECT 113.255 183.465 113.425 183.635 ;
        RECT 113.715 183.465 113.885 183.635 ;
        RECT 114.175 183.465 114.345 183.635 ;
        RECT 114.635 183.465 114.805 183.635 ;
        RECT 115.095 183.465 115.265 183.635 ;
        RECT 115.555 183.465 115.725 183.635 ;
        RECT 116.015 183.465 116.185 183.635 ;
        RECT 116.475 183.465 116.645 183.635 ;
        RECT 116.935 183.465 117.105 183.635 ;
        RECT 117.395 183.465 117.565 183.635 ;
        RECT 117.855 183.465 118.025 183.635 ;
        RECT 118.315 183.465 118.485 183.635 ;
        RECT 118.775 183.465 118.945 183.635 ;
        RECT 119.235 183.465 119.405 183.635 ;
        RECT 87.035 182.275 87.205 182.445 ;
        RECT 90.255 182.955 90.425 183.125 ;
        RECT 93.935 182.955 94.105 183.125 ;
        RECT 92.555 181.935 92.725 182.105 ;
        RECT 95.775 181.935 95.945 182.105 ;
        RECT 96.695 181.935 96.865 182.105 ;
        RECT 94.855 181.255 95.025 181.425 ;
        RECT 97.615 181.595 97.785 181.765 ;
        RECT 104.055 181.595 104.225 181.765 ;
        RECT 104.975 181.595 105.145 181.765 ;
        RECT 105.895 181.595 106.065 181.765 ;
        RECT 114.175 181.935 114.345 182.105 ;
        RECT 114.635 181.935 114.805 182.105 ;
        RECT 113.715 181.255 113.885 181.425 ;
        RECT 117.855 182.275 118.025 182.445 ;
        RECT 71.395 180.745 71.565 180.915 ;
        RECT 71.855 180.745 72.025 180.915 ;
        RECT 72.315 180.745 72.485 180.915 ;
        RECT 72.775 180.745 72.945 180.915 ;
        RECT 73.235 180.745 73.405 180.915 ;
        RECT 73.695 180.745 73.865 180.915 ;
        RECT 74.155 180.745 74.325 180.915 ;
        RECT 74.615 180.745 74.785 180.915 ;
        RECT 75.075 180.745 75.245 180.915 ;
        RECT 75.535 180.745 75.705 180.915 ;
        RECT 75.995 180.745 76.165 180.915 ;
        RECT 76.455 180.745 76.625 180.915 ;
        RECT 76.915 180.745 77.085 180.915 ;
        RECT 77.375 180.745 77.545 180.915 ;
        RECT 77.835 180.745 78.005 180.915 ;
        RECT 78.295 180.745 78.465 180.915 ;
        RECT 78.755 180.745 78.925 180.915 ;
        RECT 79.215 180.745 79.385 180.915 ;
        RECT 79.675 180.745 79.845 180.915 ;
        RECT 80.135 180.745 80.305 180.915 ;
        RECT 80.595 180.745 80.765 180.915 ;
        RECT 81.055 180.745 81.225 180.915 ;
        RECT 81.515 180.745 81.685 180.915 ;
        RECT 81.975 180.745 82.145 180.915 ;
        RECT 82.435 180.745 82.605 180.915 ;
        RECT 82.895 180.745 83.065 180.915 ;
        RECT 83.355 180.745 83.525 180.915 ;
        RECT 83.815 180.745 83.985 180.915 ;
        RECT 84.275 180.745 84.445 180.915 ;
        RECT 84.735 180.745 84.905 180.915 ;
        RECT 85.195 180.745 85.365 180.915 ;
        RECT 85.655 180.745 85.825 180.915 ;
        RECT 86.115 180.745 86.285 180.915 ;
        RECT 86.575 180.745 86.745 180.915 ;
        RECT 87.035 180.745 87.205 180.915 ;
        RECT 87.495 180.745 87.665 180.915 ;
        RECT 87.955 180.745 88.125 180.915 ;
        RECT 88.415 180.745 88.585 180.915 ;
        RECT 88.875 180.745 89.045 180.915 ;
        RECT 89.335 180.745 89.505 180.915 ;
        RECT 89.795 180.745 89.965 180.915 ;
        RECT 90.255 180.745 90.425 180.915 ;
        RECT 90.715 180.745 90.885 180.915 ;
        RECT 91.175 180.745 91.345 180.915 ;
        RECT 91.635 180.745 91.805 180.915 ;
        RECT 92.095 180.745 92.265 180.915 ;
        RECT 92.555 180.745 92.725 180.915 ;
        RECT 93.015 180.745 93.185 180.915 ;
        RECT 93.475 180.745 93.645 180.915 ;
        RECT 93.935 180.745 94.105 180.915 ;
        RECT 94.395 180.745 94.565 180.915 ;
        RECT 94.855 180.745 95.025 180.915 ;
        RECT 95.315 180.745 95.485 180.915 ;
        RECT 95.775 180.745 95.945 180.915 ;
        RECT 96.235 180.745 96.405 180.915 ;
        RECT 96.695 180.745 96.865 180.915 ;
        RECT 97.155 180.745 97.325 180.915 ;
        RECT 97.615 180.745 97.785 180.915 ;
        RECT 98.075 180.745 98.245 180.915 ;
        RECT 98.535 180.745 98.705 180.915 ;
        RECT 98.995 180.745 99.165 180.915 ;
        RECT 99.455 180.745 99.625 180.915 ;
        RECT 99.915 180.745 100.085 180.915 ;
        RECT 100.375 180.745 100.545 180.915 ;
        RECT 100.835 180.745 101.005 180.915 ;
        RECT 101.295 180.745 101.465 180.915 ;
        RECT 101.755 180.745 101.925 180.915 ;
        RECT 102.215 180.745 102.385 180.915 ;
        RECT 102.675 180.745 102.845 180.915 ;
        RECT 103.135 180.745 103.305 180.915 ;
        RECT 103.595 180.745 103.765 180.915 ;
        RECT 104.055 180.745 104.225 180.915 ;
        RECT 104.515 180.745 104.685 180.915 ;
        RECT 104.975 180.745 105.145 180.915 ;
        RECT 105.435 180.745 105.605 180.915 ;
        RECT 105.895 180.745 106.065 180.915 ;
        RECT 106.355 180.745 106.525 180.915 ;
        RECT 106.815 180.745 106.985 180.915 ;
        RECT 107.275 180.745 107.445 180.915 ;
        RECT 107.735 180.745 107.905 180.915 ;
        RECT 108.195 180.745 108.365 180.915 ;
        RECT 108.655 180.745 108.825 180.915 ;
        RECT 109.115 180.745 109.285 180.915 ;
        RECT 109.575 180.745 109.745 180.915 ;
        RECT 110.035 180.745 110.205 180.915 ;
        RECT 110.495 180.745 110.665 180.915 ;
        RECT 110.955 180.745 111.125 180.915 ;
        RECT 111.415 180.745 111.585 180.915 ;
        RECT 111.875 180.745 112.045 180.915 ;
        RECT 112.335 180.745 112.505 180.915 ;
        RECT 112.795 180.745 112.965 180.915 ;
        RECT 113.255 180.745 113.425 180.915 ;
        RECT 113.715 180.745 113.885 180.915 ;
        RECT 114.175 180.745 114.345 180.915 ;
        RECT 114.635 180.745 114.805 180.915 ;
        RECT 115.095 180.745 115.265 180.915 ;
        RECT 115.555 180.745 115.725 180.915 ;
        RECT 116.015 180.745 116.185 180.915 ;
        RECT 116.475 180.745 116.645 180.915 ;
        RECT 116.935 180.745 117.105 180.915 ;
        RECT 117.395 180.745 117.565 180.915 ;
        RECT 117.855 180.745 118.025 180.915 ;
        RECT 118.315 180.745 118.485 180.915 ;
        RECT 118.775 180.745 118.945 180.915 ;
        RECT 119.235 180.745 119.405 180.915 ;
        RECT 73.695 179.555 73.865 179.725 ;
        RECT 74.160 179.555 74.330 179.725 ;
        RECT 75.075 179.215 75.245 179.385 ;
        RECT 74.565 178.875 74.735 179.045 ;
        RECT 75.995 179.555 76.165 179.725 ;
        RECT 77.355 179.895 77.525 180.065 ;
        RECT 77.715 179.895 77.885 180.065 ;
        RECT 76.455 178.875 76.625 179.045 ;
        RECT 79.575 179.555 79.745 179.725 ;
        RECT 80.955 179.895 81.125 180.065 ;
        RECT 80.655 179.580 80.825 179.750 ;
        RECT 79.575 178.875 79.745 179.045 ;
        RECT 82.435 178.875 82.605 179.045 ;
        RECT 86.115 179.555 86.285 179.725 ;
        RECT 85.195 178.535 85.365 178.705 ;
        RECT 98.535 179.895 98.705 180.065 ;
        RECT 99.455 179.555 99.625 179.725 ;
        RECT 101.295 180.235 101.465 180.405 ;
        RECT 97.615 178.535 97.785 178.705 ;
        RECT 102.215 179.555 102.385 179.725 ;
        RECT 103.135 179.555 103.305 179.725 ;
        RECT 103.595 179.555 103.765 179.725 ;
        RECT 105.435 179.555 105.605 179.725 ;
        RECT 105.920 178.875 106.090 179.045 ;
        RECT 106.315 179.215 106.485 179.385 ;
        RECT 106.770 179.555 106.940 179.725 ;
        RECT 107.505 179.215 107.675 179.385 ;
        RECT 108.020 178.875 108.190 179.045 ;
        RECT 109.590 178.875 109.760 179.045 ;
        RECT 110.025 179.215 110.195 179.385 ;
        RECT 112.335 178.535 112.505 178.705 ;
        RECT 71.395 178.025 71.565 178.195 ;
        RECT 71.855 178.025 72.025 178.195 ;
        RECT 72.315 178.025 72.485 178.195 ;
        RECT 72.775 178.025 72.945 178.195 ;
        RECT 73.235 178.025 73.405 178.195 ;
        RECT 73.695 178.025 73.865 178.195 ;
        RECT 74.155 178.025 74.325 178.195 ;
        RECT 74.615 178.025 74.785 178.195 ;
        RECT 75.075 178.025 75.245 178.195 ;
        RECT 75.535 178.025 75.705 178.195 ;
        RECT 75.995 178.025 76.165 178.195 ;
        RECT 76.455 178.025 76.625 178.195 ;
        RECT 76.915 178.025 77.085 178.195 ;
        RECT 77.375 178.025 77.545 178.195 ;
        RECT 77.835 178.025 78.005 178.195 ;
        RECT 78.295 178.025 78.465 178.195 ;
        RECT 78.755 178.025 78.925 178.195 ;
        RECT 79.215 178.025 79.385 178.195 ;
        RECT 79.675 178.025 79.845 178.195 ;
        RECT 80.135 178.025 80.305 178.195 ;
        RECT 80.595 178.025 80.765 178.195 ;
        RECT 81.055 178.025 81.225 178.195 ;
        RECT 81.515 178.025 81.685 178.195 ;
        RECT 81.975 178.025 82.145 178.195 ;
        RECT 82.435 178.025 82.605 178.195 ;
        RECT 82.895 178.025 83.065 178.195 ;
        RECT 83.355 178.025 83.525 178.195 ;
        RECT 83.815 178.025 83.985 178.195 ;
        RECT 84.275 178.025 84.445 178.195 ;
        RECT 84.735 178.025 84.905 178.195 ;
        RECT 85.195 178.025 85.365 178.195 ;
        RECT 85.655 178.025 85.825 178.195 ;
        RECT 86.115 178.025 86.285 178.195 ;
        RECT 86.575 178.025 86.745 178.195 ;
        RECT 87.035 178.025 87.205 178.195 ;
        RECT 87.495 178.025 87.665 178.195 ;
        RECT 87.955 178.025 88.125 178.195 ;
        RECT 88.415 178.025 88.585 178.195 ;
        RECT 88.875 178.025 89.045 178.195 ;
        RECT 89.335 178.025 89.505 178.195 ;
        RECT 89.795 178.025 89.965 178.195 ;
        RECT 90.255 178.025 90.425 178.195 ;
        RECT 90.715 178.025 90.885 178.195 ;
        RECT 91.175 178.025 91.345 178.195 ;
        RECT 91.635 178.025 91.805 178.195 ;
        RECT 92.095 178.025 92.265 178.195 ;
        RECT 92.555 178.025 92.725 178.195 ;
        RECT 93.015 178.025 93.185 178.195 ;
        RECT 93.475 178.025 93.645 178.195 ;
        RECT 93.935 178.025 94.105 178.195 ;
        RECT 94.395 178.025 94.565 178.195 ;
        RECT 94.855 178.025 95.025 178.195 ;
        RECT 95.315 178.025 95.485 178.195 ;
        RECT 95.775 178.025 95.945 178.195 ;
        RECT 96.235 178.025 96.405 178.195 ;
        RECT 96.695 178.025 96.865 178.195 ;
        RECT 97.155 178.025 97.325 178.195 ;
        RECT 97.615 178.025 97.785 178.195 ;
        RECT 98.075 178.025 98.245 178.195 ;
        RECT 98.535 178.025 98.705 178.195 ;
        RECT 98.995 178.025 99.165 178.195 ;
        RECT 99.455 178.025 99.625 178.195 ;
        RECT 99.915 178.025 100.085 178.195 ;
        RECT 100.375 178.025 100.545 178.195 ;
        RECT 100.835 178.025 101.005 178.195 ;
        RECT 101.295 178.025 101.465 178.195 ;
        RECT 101.755 178.025 101.925 178.195 ;
        RECT 102.215 178.025 102.385 178.195 ;
        RECT 102.675 178.025 102.845 178.195 ;
        RECT 103.135 178.025 103.305 178.195 ;
        RECT 103.595 178.025 103.765 178.195 ;
        RECT 104.055 178.025 104.225 178.195 ;
        RECT 104.515 178.025 104.685 178.195 ;
        RECT 104.975 178.025 105.145 178.195 ;
        RECT 105.435 178.025 105.605 178.195 ;
        RECT 105.895 178.025 106.065 178.195 ;
        RECT 106.355 178.025 106.525 178.195 ;
        RECT 106.815 178.025 106.985 178.195 ;
        RECT 107.275 178.025 107.445 178.195 ;
        RECT 107.735 178.025 107.905 178.195 ;
        RECT 108.195 178.025 108.365 178.195 ;
        RECT 108.655 178.025 108.825 178.195 ;
        RECT 109.115 178.025 109.285 178.195 ;
        RECT 109.575 178.025 109.745 178.195 ;
        RECT 110.035 178.025 110.205 178.195 ;
        RECT 110.495 178.025 110.665 178.195 ;
        RECT 110.955 178.025 111.125 178.195 ;
        RECT 111.415 178.025 111.585 178.195 ;
        RECT 111.875 178.025 112.045 178.195 ;
        RECT 112.335 178.025 112.505 178.195 ;
        RECT 112.795 178.025 112.965 178.195 ;
        RECT 113.255 178.025 113.425 178.195 ;
        RECT 113.715 178.025 113.885 178.195 ;
        RECT 114.175 178.025 114.345 178.195 ;
        RECT 114.635 178.025 114.805 178.195 ;
        RECT 115.095 178.025 115.265 178.195 ;
        RECT 115.555 178.025 115.725 178.195 ;
        RECT 116.015 178.025 116.185 178.195 ;
        RECT 116.475 178.025 116.645 178.195 ;
        RECT 116.935 178.025 117.105 178.195 ;
        RECT 117.395 178.025 117.565 178.195 ;
        RECT 117.855 178.025 118.025 178.195 ;
        RECT 118.315 178.025 118.485 178.195 ;
        RECT 118.775 178.025 118.945 178.195 ;
        RECT 119.235 178.025 119.405 178.195 ;
        RECT 73.695 177.515 73.865 177.685 ;
        RECT 75.075 176.835 75.245 177.005 ;
        RECT 75.535 176.495 75.705 176.665 ;
        RECT 81.055 176.835 81.225 177.005 ;
        RECT 83.355 176.835 83.525 177.005 ;
        RECT 82.895 176.495 83.065 176.665 ;
        RECT 99.455 177.515 99.625 177.685 ;
        RECT 101.295 177.515 101.465 177.685 ;
        RECT 92.095 176.155 92.265 176.325 ;
        RECT 104.055 176.495 104.225 176.665 ;
        RECT 105.435 175.815 105.605 175.985 ;
        RECT 108.655 176.495 108.825 176.665 ;
        RECT 110.495 175.815 110.665 175.985 ;
        RECT 113.255 176.835 113.425 177.005 ;
        RECT 115.095 177.515 115.265 177.685 ;
        RECT 114.635 176.495 114.805 176.665 ;
        RECT 112.795 175.815 112.965 175.985 ;
        RECT 115.555 176.495 115.725 176.665 ;
        RECT 116.015 176.495 116.185 176.665 ;
        RECT 116.935 176.495 117.105 176.665 ;
        RECT 116.015 175.815 116.185 175.985 ;
        RECT 71.395 175.305 71.565 175.475 ;
        RECT 71.855 175.305 72.025 175.475 ;
        RECT 72.315 175.305 72.485 175.475 ;
        RECT 72.775 175.305 72.945 175.475 ;
        RECT 73.235 175.305 73.405 175.475 ;
        RECT 73.695 175.305 73.865 175.475 ;
        RECT 74.155 175.305 74.325 175.475 ;
        RECT 74.615 175.305 74.785 175.475 ;
        RECT 75.075 175.305 75.245 175.475 ;
        RECT 75.535 175.305 75.705 175.475 ;
        RECT 75.995 175.305 76.165 175.475 ;
        RECT 76.455 175.305 76.625 175.475 ;
        RECT 76.915 175.305 77.085 175.475 ;
        RECT 77.375 175.305 77.545 175.475 ;
        RECT 77.835 175.305 78.005 175.475 ;
        RECT 78.295 175.305 78.465 175.475 ;
        RECT 78.755 175.305 78.925 175.475 ;
        RECT 79.215 175.305 79.385 175.475 ;
        RECT 79.675 175.305 79.845 175.475 ;
        RECT 80.135 175.305 80.305 175.475 ;
        RECT 80.595 175.305 80.765 175.475 ;
        RECT 81.055 175.305 81.225 175.475 ;
        RECT 81.515 175.305 81.685 175.475 ;
        RECT 81.975 175.305 82.145 175.475 ;
        RECT 82.435 175.305 82.605 175.475 ;
        RECT 82.895 175.305 83.065 175.475 ;
        RECT 83.355 175.305 83.525 175.475 ;
        RECT 83.815 175.305 83.985 175.475 ;
        RECT 84.275 175.305 84.445 175.475 ;
        RECT 84.735 175.305 84.905 175.475 ;
        RECT 85.195 175.305 85.365 175.475 ;
        RECT 85.655 175.305 85.825 175.475 ;
        RECT 86.115 175.305 86.285 175.475 ;
        RECT 86.575 175.305 86.745 175.475 ;
        RECT 87.035 175.305 87.205 175.475 ;
        RECT 87.495 175.305 87.665 175.475 ;
        RECT 87.955 175.305 88.125 175.475 ;
        RECT 88.415 175.305 88.585 175.475 ;
        RECT 88.875 175.305 89.045 175.475 ;
        RECT 89.335 175.305 89.505 175.475 ;
        RECT 89.795 175.305 89.965 175.475 ;
        RECT 90.255 175.305 90.425 175.475 ;
        RECT 90.715 175.305 90.885 175.475 ;
        RECT 91.175 175.305 91.345 175.475 ;
        RECT 91.635 175.305 91.805 175.475 ;
        RECT 92.095 175.305 92.265 175.475 ;
        RECT 92.555 175.305 92.725 175.475 ;
        RECT 93.015 175.305 93.185 175.475 ;
        RECT 93.475 175.305 93.645 175.475 ;
        RECT 93.935 175.305 94.105 175.475 ;
        RECT 94.395 175.305 94.565 175.475 ;
        RECT 94.855 175.305 95.025 175.475 ;
        RECT 95.315 175.305 95.485 175.475 ;
        RECT 95.775 175.305 95.945 175.475 ;
        RECT 96.235 175.305 96.405 175.475 ;
        RECT 96.695 175.305 96.865 175.475 ;
        RECT 97.155 175.305 97.325 175.475 ;
        RECT 97.615 175.305 97.785 175.475 ;
        RECT 98.075 175.305 98.245 175.475 ;
        RECT 98.535 175.305 98.705 175.475 ;
        RECT 98.995 175.305 99.165 175.475 ;
        RECT 99.455 175.305 99.625 175.475 ;
        RECT 99.915 175.305 100.085 175.475 ;
        RECT 100.375 175.305 100.545 175.475 ;
        RECT 100.835 175.305 101.005 175.475 ;
        RECT 101.295 175.305 101.465 175.475 ;
        RECT 101.755 175.305 101.925 175.475 ;
        RECT 102.215 175.305 102.385 175.475 ;
        RECT 102.675 175.305 102.845 175.475 ;
        RECT 103.135 175.305 103.305 175.475 ;
        RECT 103.595 175.305 103.765 175.475 ;
        RECT 104.055 175.305 104.225 175.475 ;
        RECT 104.515 175.305 104.685 175.475 ;
        RECT 104.975 175.305 105.145 175.475 ;
        RECT 105.435 175.305 105.605 175.475 ;
        RECT 105.895 175.305 106.065 175.475 ;
        RECT 106.355 175.305 106.525 175.475 ;
        RECT 106.815 175.305 106.985 175.475 ;
        RECT 107.275 175.305 107.445 175.475 ;
        RECT 107.735 175.305 107.905 175.475 ;
        RECT 108.195 175.305 108.365 175.475 ;
        RECT 108.655 175.305 108.825 175.475 ;
        RECT 109.115 175.305 109.285 175.475 ;
        RECT 109.575 175.305 109.745 175.475 ;
        RECT 110.035 175.305 110.205 175.475 ;
        RECT 110.495 175.305 110.665 175.475 ;
        RECT 110.955 175.305 111.125 175.475 ;
        RECT 111.415 175.305 111.585 175.475 ;
        RECT 111.875 175.305 112.045 175.475 ;
        RECT 112.335 175.305 112.505 175.475 ;
        RECT 112.795 175.305 112.965 175.475 ;
        RECT 113.255 175.305 113.425 175.475 ;
        RECT 113.715 175.305 113.885 175.475 ;
        RECT 114.175 175.305 114.345 175.475 ;
        RECT 114.635 175.305 114.805 175.475 ;
        RECT 115.095 175.305 115.265 175.475 ;
        RECT 115.555 175.305 115.725 175.475 ;
        RECT 116.015 175.305 116.185 175.475 ;
        RECT 116.475 175.305 116.645 175.475 ;
        RECT 116.935 175.305 117.105 175.475 ;
        RECT 117.395 175.305 117.565 175.475 ;
        RECT 117.855 175.305 118.025 175.475 ;
        RECT 118.315 175.305 118.485 175.475 ;
        RECT 118.775 175.305 118.945 175.475 ;
        RECT 119.235 175.305 119.405 175.475 ;
        RECT 74.155 174.115 74.325 174.285 ;
        RECT 74.620 174.115 74.790 174.285 ;
        RECT 75.535 173.775 75.705 173.945 ;
        RECT 75.025 173.435 75.195 173.605 ;
        RECT 76.455 174.115 76.625 174.285 ;
        RECT 77.815 174.455 77.985 174.625 ;
        RECT 78.175 174.455 78.345 174.625 ;
        RECT 76.915 173.435 77.085 173.605 ;
        RECT 80.035 174.115 80.205 174.285 ;
        RECT 81.415 174.455 81.585 174.625 ;
        RECT 81.115 174.140 81.285 174.310 ;
        RECT 80.035 173.435 80.205 173.605 ;
        RECT 82.895 173.095 83.065 173.265 ;
        RECT 84.735 174.115 84.905 174.285 ;
        RECT 85.200 174.115 85.370 174.285 ;
        RECT 86.115 173.775 86.285 173.945 ;
        RECT 85.605 173.435 85.775 173.605 ;
        RECT 87.035 174.115 87.205 174.285 ;
        RECT 88.395 174.455 88.565 174.625 ;
        RECT 88.755 174.455 88.925 174.625 ;
        RECT 87.495 173.435 87.665 173.605 ;
        RECT 90.615 174.115 90.785 174.285 ;
        RECT 91.995 174.455 92.165 174.625 ;
        RECT 91.695 174.140 91.865 174.310 ;
        RECT 90.615 173.435 90.785 173.605 ;
        RECT 93.475 173.095 93.645 173.265 ;
        RECT 95.315 174.115 95.485 174.285 ;
        RECT 94.395 173.435 94.565 173.605 ;
        RECT 97.615 174.115 97.785 174.285 ;
        RECT 96.235 173.095 96.405 173.265 ;
        RECT 98.100 173.435 98.270 173.605 ;
        RECT 98.495 173.775 98.665 173.945 ;
        RECT 98.895 174.115 99.065 174.285 ;
        RECT 99.685 173.775 99.855 173.945 ;
        RECT 100.200 173.435 100.370 173.605 ;
        RECT 101.770 173.435 101.940 173.605 ;
        RECT 102.205 173.775 102.375 173.945 ;
        RECT 104.515 174.795 104.685 174.965 ;
        RECT 106.355 173.775 106.525 173.945 ;
        RECT 107.275 174.795 107.445 174.965 ;
        RECT 109.115 174.795 109.285 174.965 ;
        RECT 106.815 173.775 106.985 173.945 ;
        RECT 109.575 174.115 109.745 174.285 ;
        RECT 112.795 174.455 112.965 174.625 ;
        RECT 110.495 174.115 110.665 174.285 ;
        RECT 110.495 173.095 110.665 173.265 ;
        RECT 111.875 173.775 112.045 173.945 ;
        RECT 113.255 174.795 113.425 174.965 ;
        RECT 115.095 173.095 115.265 173.265 ;
        RECT 116.475 174.455 116.645 174.625 ;
        RECT 117.395 174.115 117.565 174.285 ;
        RECT 115.555 173.095 115.725 173.265 ;
        RECT 71.395 172.585 71.565 172.755 ;
        RECT 71.855 172.585 72.025 172.755 ;
        RECT 72.315 172.585 72.485 172.755 ;
        RECT 72.775 172.585 72.945 172.755 ;
        RECT 73.235 172.585 73.405 172.755 ;
        RECT 73.695 172.585 73.865 172.755 ;
        RECT 74.155 172.585 74.325 172.755 ;
        RECT 74.615 172.585 74.785 172.755 ;
        RECT 75.075 172.585 75.245 172.755 ;
        RECT 75.535 172.585 75.705 172.755 ;
        RECT 75.995 172.585 76.165 172.755 ;
        RECT 76.455 172.585 76.625 172.755 ;
        RECT 76.915 172.585 77.085 172.755 ;
        RECT 77.375 172.585 77.545 172.755 ;
        RECT 77.835 172.585 78.005 172.755 ;
        RECT 78.295 172.585 78.465 172.755 ;
        RECT 78.755 172.585 78.925 172.755 ;
        RECT 79.215 172.585 79.385 172.755 ;
        RECT 79.675 172.585 79.845 172.755 ;
        RECT 80.135 172.585 80.305 172.755 ;
        RECT 80.595 172.585 80.765 172.755 ;
        RECT 81.055 172.585 81.225 172.755 ;
        RECT 81.515 172.585 81.685 172.755 ;
        RECT 81.975 172.585 82.145 172.755 ;
        RECT 82.435 172.585 82.605 172.755 ;
        RECT 82.895 172.585 83.065 172.755 ;
        RECT 83.355 172.585 83.525 172.755 ;
        RECT 83.815 172.585 83.985 172.755 ;
        RECT 84.275 172.585 84.445 172.755 ;
        RECT 84.735 172.585 84.905 172.755 ;
        RECT 85.195 172.585 85.365 172.755 ;
        RECT 85.655 172.585 85.825 172.755 ;
        RECT 86.115 172.585 86.285 172.755 ;
        RECT 86.575 172.585 86.745 172.755 ;
        RECT 87.035 172.585 87.205 172.755 ;
        RECT 87.495 172.585 87.665 172.755 ;
        RECT 87.955 172.585 88.125 172.755 ;
        RECT 88.415 172.585 88.585 172.755 ;
        RECT 88.875 172.585 89.045 172.755 ;
        RECT 89.335 172.585 89.505 172.755 ;
        RECT 89.795 172.585 89.965 172.755 ;
        RECT 90.255 172.585 90.425 172.755 ;
        RECT 90.715 172.585 90.885 172.755 ;
        RECT 91.175 172.585 91.345 172.755 ;
        RECT 91.635 172.585 91.805 172.755 ;
        RECT 92.095 172.585 92.265 172.755 ;
        RECT 92.555 172.585 92.725 172.755 ;
        RECT 93.015 172.585 93.185 172.755 ;
        RECT 93.475 172.585 93.645 172.755 ;
        RECT 93.935 172.585 94.105 172.755 ;
        RECT 94.395 172.585 94.565 172.755 ;
        RECT 94.855 172.585 95.025 172.755 ;
        RECT 95.315 172.585 95.485 172.755 ;
        RECT 95.775 172.585 95.945 172.755 ;
        RECT 96.235 172.585 96.405 172.755 ;
        RECT 96.695 172.585 96.865 172.755 ;
        RECT 97.155 172.585 97.325 172.755 ;
        RECT 97.615 172.585 97.785 172.755 ;
        RECT 98.075 172.585 98.245 172.755 ;
        RECT 98.535 172.585 98.705 172.755 ;
        RECT 98.995 172.585 99.165 172.755 ;
        RECT 99.455 172.585 99.625 172.755 ;
        RECT 99.915 172.585 100.085 172.755 ;
        RECT 100.375 172.585 100.545 172.755 ;
        RECT 100.835 172.585 101.005 172.755 ;
        RECT 101.295 172.585 101.465 172.755 ;
        RECT 101.755 172.585 101.925 172.755 ;
        RECT 102.215 172.585 102.385 172.755 ;
        RECT 102.675 172.585 102.845 172.755 ;
        RECT 103.135 172.585 103.305 172.755 ;
        RECT 103.595 172.585 103.765 172.755 ;
        RECT 104.055 172.585 104.225 172.755 ;
        RECT 104.515 172.585 104.685 172.755 ;
        RECT 104.975 172.585 105.145 172.755 ;
        RECT 105.435 172.585 105.605 172.755 ;
        RECT 105.895 172.585 106.065 172.755 ;
        RECT 106.355 172.585 106.525 172.755 ;
        RECT 106.815 172.585 106.985 172.755 ;
        RECT 107.275 172.585 107.445 172.755 ;
        RECT 107.735 172.585 107.905 172.755 ;
        RECT 108.195 172.585 108.365 172.755 ;
        RECT 108.655 172.585 108.825 172.755 ;
        RECT 109.115 172.585 109.285 172.755 ;
        RECT 109.575 172.585 109.745 172.755 ;
        RECT 110.035 172.585 110.205 172.755 ;
        RECT 110.495 172.585 110.665 172.755 ;
        RECT 110.955 172.585 111.125 172.755 ;
        RECT 111.415 172.585 111.585 172.755 ;
        RECT 111.875 172.585 112.045 172.755 ;
        RECT 112.335 172.585 112.505 172.755 ;
        RECT 112.795 172.585 112.965 172.755 ;
        RECT 113.255 172.585 113.425 172.755 ;
        RECT 113.715 172.585 113.885 172.755 ;
        RECT 114.175 172.585 114.345 172.755 ;
        RECT 114.635 172.585 114.805 172.755 ;
        RECT 115.095 172.585 115.265 172.755 ;
        RECT 115.555 172.585 115.725 172.755 ;
        RECT 116.015 172.585 116.185 172.755 ;
        RECT 116.475 172.585 116.645 172.755 ;
        RECT 116.935 172.585 117.105 172.755 ;
        RECT 117.395 172.585 117.565 172.755 ;
        RECT 117.855 172.585 118.025 172.755 ;
        RECT 118.315 172.585 118.485 172.755 ;
        RECT 118.775 172.585 118.945 172.755 ;
        RECT 119.235 172.585 119.405 172.755 ;
        RECT 75.535 172.075 75.705 172.245 ;
        RECT 76.455 171.395 76.625 171.565 ;
        RECT 76.915 171.055 77.085 171.225 ;
        RECT 85.655 172.075 85.825 172.245 ;
        RECT 84.735 171.055 84.905 171.225 ;
        RECT 90.715 171.395 90.885 171.565 ;
        RECT 92.095 171.395 92.265 171.565 ;
        RECT 103.160 171.735 103.330 171.905 ;
        RECT 92.555 170.715 92.725 170.885 ;
        RECT 102.675 171.055 102.845 171.225 ;
        RECT 98.995 170.375 99.165 170.545 ;
        RECT 103.555 171.395 103.725 171.565 ;
        RECT 103.900 170.715 104.070 170.885 ;
        RECT 105.260 171.735 105.430 171.905 ;
        RECT 104.745 171.395 104.915 171.565 ;
        RECT 106.830 171.735 107.000 171.905 ;
        RECT 107.265 171.395 107.435 171.565 ;
        RECT 109.575 171.735 109.745 171.905 ;
        RECT 110.495 172.075 110.665 172.245 ;
        RECT 113.255 171.395 113.425 171.565 ;
        RECT 114.175 170.375 114.345 170.545 ;
        RECT 116.935 171.395 117.105 171.565 ;
        RECT 71.395 169.865 71.565 170.035 ;
        RECT 71.855 169.865 72.025 170.035 ;
        RECT 72.315 169.865 72.485 170.035 ;
        RECT 72.775 169.865 72.945 170.035 ;
        RECT 73.235 169.865 73.405 170.035 ;
        RECT 73.695 169.865 73.865 170.035 ;
        RECT 74.155 169.865 74.325 170.035 ;
        RECT 74.615 169.865 74.785 170.035 ;
        RECT 75.075 169.865 75.245 170.035 ;
        RECT 75.535 169.865 75.705 170.035 ;
        RECT 75.995 169.865 76.165 170.035 ;
        RECT 76.455 169.865 76.625 170.035 ;
        RECT 76.915 169.865 77.085 170.035 ;
        RECT 77.375 169.865 77.545 170.035 ;
        RECT 77.835 169.865 78.005 170.035 ;
        RECT 78.295 169.865 78.465 170.035 ;
        RECT 78.755 169.865 78.925 170.035 ;
        RECT 79.215 169.865 79.385 170.035 ;
        RECT 79.675 169.865 79.845 170.035 ;
        RECT 80.135 169.865 80.305 170.035 ;
        RECT 80.595 169.865 80.765 170.035 ;
        RECT 81.055 169.865 81.225 170.035 ;
        RECT 81.515 169.865 81.685 170.035 ;
        RECT 81.975 169.865 82.145 170.035 ;
        RECT 82.435 169.865 82.605 170.035 ;
        RECT 82.895 169.865 83.065 170.035 ;
        RECT 83.355 169.865 83.525 170.035 ;
        RECT 83.815 169.865 83.985 170.035 ;
        RECT 84.275 169.865 84.445 170.035 ;
        RECT 84.735 169.865 84.905 170.035 ;
        RECT 85.195 169.865 85.365 170.035 ;
        RECT 85.655 169.865 85.825 170.035 ;
        RECT 86.115 169.865 86.285 170.035 ;
        RECT 86.575 169.865 86.745 170.035 ;
        RECT 87.035 169.865 87.205 170.035 ;
        RECT 87.495 169.865 87.665 170.035 ;
        RECT 87.955 169.865 88.125 170.035 ;
        RECT 88.415 169.865 88.585 170.035 ;
        RECT 88.875 169.865 89.045 170.035 ;
        RECT 89.335 169.865 89.505 170.035 ;
        RECT 89.795 169.865 89.965 170.035 ;
        RECT 90.255 169.865 90.425 170.035 ;
        RECT 90.715 169.865 90.885 170.035 ;
        RECT 91.175 169.865 91.345 170.035 ;
        RECT 91.635 169.865 91.805 170.035 ;
        RECT 92.095 169.865 92.265 170.035 ;
        RECT 92.555 169.865 92.725 170.035 ;
        RECT 93.015 169.865 93.185 170.035 ;
        RECT 93.475 169.865 93.645 170.035 ;
        RECT 93.935 169.865 94.105 170.035 ;
        RECT 94.395 169.865 94.565 170.035 ;
        RECT 94.855 169.865 95.025 170.035 ;
        RECT 95.315 169.865 95.485 170.035 ;
        RECT 95.775 169.865 95.945 170.035 ;
        RECT 96.235 169.865 96.405 170.035 ;
        RECT 96.695 169.865 96.865 170.035 ;
        RECT 97.155 169.865 97.325 170.035 ;
        RECT 97.615 169.865 97.785 170.035 ;
        RECT 98.075 169.865 98.245 170.035 ;
        RECT 98.535 169.865 98.705 170.035 ;
        RECT 98.995 169.865 99.165 170.035 ;
        RECT 99.455 169.865 99.625 170.035 ;
        RECT 99.915 169.865 100.085 170.035 ;
        RECT 100.375 169.865 100.545 170.035 ;
        RECT 100.835 169.865 101.005 170.035 ;
        RECT 101.295 169.865 101.465 170.035 ;
        RECT 101.755 169.865 101.925 170.035 ;
        RECT 102.215 169.865 102.385 170.035 ;
        RECT 102.675 169.865 102.845 170.035 ;
        RECT 103.135 169.865 103.305 170.035 ;
        RECT 103.595 169.865 103.765 170.035 ;
        RECT 104.055 169.865 104.225 170.035 ;
        RECT 104.515 169.865 104.685 170.035 ;
        RECT 104.975 169.865 105.145 170.035 ;
        RECT 105.435 169.865 105.605 170.035 ;
        RECT 105.895 169.865 106.065 170.035 ;
        RECT 106.355 169.865 106.525 170.035 ;
        RECT 106.815 169.865 106.985 170.035 ;
        RECT 107.275 169.865 107.445 170.035 ;
        RECT 107.735 169.865 107.905 170.035 ;
        RECT 108.195 169.865 108.365 170.035 ;
        RECT 108.655 169.865 108.825 170.035 ;
        RECT 109.115 169.865 109.285 170.035 ;
        RECT 109.575 169.865 109.745 170.035 ;
        RECT 110.035 169.865 110.205 170.035 ;
        RECT 110.495 169.865 110.665 170.035 ;
        RECT 110.955 169.865 111.125 170.035 ;
        RECT 111.415 169.865 111.585 170.035 ;
        RECT 111.875 169.865 112.045 170.035 ;
        RECT 112.335 169.865 112.505 170.035 ;
        RECT 112.795 169.865 112.965 170.035 ;
        RECT 113.255 169.865 113.425 170.035 ;
        RECT 113.715 169.865 113.885 170.035 ;
        RECT 114.175 169.865 114.345 170.035 ;
        RECT 114.635 169.865 114.805 170.035 ;
        RECT 115.095 169.865 115.265 170.035 ;
        RECT 115.555 169.865 115.725 170.035 ;
        RECT 116.015 169.865 116.185 170.035 ;
        RECT 116.475 169.865 116.645 170.035 ;
        RECT 116.935 169.865 117.105 170.035 ;
        RECT 117.395 169.865 117.565 170.035 ;
        RECT 117.855 169.865 118.025 170.035 ;
        RECT 118.315 169.865 118.485 170.035 ;
        RECT 118.775 169.865 118.945 170.035 ;
        RECT 119.235 169.865 119.405 170.035 ;
        RECT 85.655 168.675 85.825 168.845 ;
        RECT 85.195 168.335 85.365 168.505 ;
        RECT 87.495 167.995 87.665 168.165 ;
        RECT 88.875 168.675 89.045 168.845 ;
        RECT 88.415 168.335 88.585 168.505 ;
        RECT 91.175 168.335 91.345 168.505 ;
        RECT 90.715 167.655 90.885 167.825 ;
        RECT 97.615 168.675 97.785 168.845 ;
        RECT 94.395 167.655 94.565 167.825 ;
        RECT 104.515 169.355 104.685 169.525 ;
        RECT 98.535 167.655 98.705 167.825 ;
        RECT 105.435 168.675 105.605 168.845 ;
        RECT 110.495 169.355 110.665 169.525 ;
        RECT 108.655 168.675 108.825 168.845 ;
        RECT 109.115 168.335 109.285 168.505 ;
        RECT 110.955 168.335 111.125 168.505 ;
        RECT 111.440 167.995 111.610 168.165 ;
        RECT 111.835 168.335 112.005 168.505 ;
        RECT 112.180 169.015 112.350 169.185 ;
        RECT 113.025 168.335 113.195 168.505 ;
        RECT 113.540 167.995 113.710 168.165 ;
        RECT 115.110 167.995 115.280 168.165 ;
        RECT 115.545 168.335 115.715 168.505 ;
        RECT 117.855 169.355 118.025 169.525 ;
        RECT 71.395 167.145 71.565 167.315 ;
        RECT 71.855 167.145 72.025 167.315 ;
        RECT 72.315 167.145 72.485 167.315 ;
        RECT 72.775 167.145 72.945 167.315 ;
        RECT 73.235 167.145 73.405 167.315 ;
        RECT 73.695 167.145 73.865 167.315 ;
        RECT 74.155 167.145 74.325 167.315 ;
        RECT 74.615 167.145 74.785 167.315 ;
        RECT 75.075 167.145 75.245 167.315 ;
        RECT 75.535 167.145 75.705 167.315 ;
        RECT 75.995 167.145 76.165 167.315 ;
        RECT 76.455 167.145 76.625 167.315 ;
        RECT 76.915 167.145 77.085 167.315 ;
        RECT 77.375 167.145 77.545 167.315 ;
        RECT 77.835 167.145 78.005 167.315 ;
        RECT 78.295 167.145 78.465 167.315 ;
        RECT 78.755 167.145 78.925 167.315 ;
        RECT 79.215 167.145 79.385 167.315 ;
        RECT 79.675 167.145 79.845 167.315 ;
        RECT 80.135 167.145 80.305 167.315 ;
        RECT 80.595 167.145 80.765 167.315 ;
        RECT 81.055 167.145 81.225 167.315 ;
        RECT 81.515 167.145 81.685 167.315 ;
        RECT 81.975 167.145 82.145 167.315 ;
        RECT 82.435 167.145 82.605 167.315 ;
        RECT 82.895 167.145 83.065 167.315 ;
        RECT 83.355 167.145 83.525 167.315 ;
        RECT 83.815 167.145 83.985 167.315 ;
        RECT 84.275 167.145 84.445 167.315 ;
        RECT 84.735 167.145 84.905 167.315 ;
        RECT 85.195 167.145 85.365 167.315 ;
        RECT 85.655 167.145 85.825 167.315 ;
        RECT 86.115 167.145 86.285 167.315 ;
        RECT 86.575 167.145 86.745 167.315 ;
        RECT 87.035 167.145 87.205 167.315 ;
        RECT 87.495 167.145 87.665 167.315 ;
        RECT 87.955 167.145 88.125 167.315 ;
        RECT 88.415 167.145 88.585 167.315 ;
        RECT 88.875 167.145 89.045 167.315 ;
        RECT 89.335 167.145 89.505 167.315 ;
        RECT 89.795 167.145 89.965 167.315 ;
        RECT 90.255 167.145 90.425 167.315 ;
        RECT 90.715 167.145 90.885 167.315 ;
        RECT 91.175 167.145 91.345 167.315 ;
        RECT 91.635 167.145 91.805 167.315 ;
        RECT 92.095 167.145 92.265 167.315 ;
        RECT 92.555 167.145 92.725 167.315 ;
        RECT 93.015 167.145 93.185 167.315 ;
        RECT 93.475 167.145 93.645 167.315 ;
        RECT 93.935 167.145 94.105 167.315 ;
        RECT 94.395 167.145 94.565 167.315 ;
        RECT 94.855 167.145 95.025 167.315 ;
        RECT 95.315 167.145 95.485 167.315 ;
        RECT 95.775 167.145 95.945 167.315 ;
        RECT 96.235 167.145 96.405 167.315 ;
        RECT 96.695 167.145 96.865 167.315 ;
        RECT 97.155 167.145 97.325 167.315 ;
        RECT 97.615 167.145 97.785 167.315 ;
        RECT 98.075 167.145 98.245 167.315 ;
        RECT 98.535 167.145 98.705 167.315 ;
        RECT 98.995 167.145 99.165 167.315 ;
        RECT 99.455 167.145 99.625 167.315 ;
        RECT 99.915 167.145 100.085 167.315 ;
        RECT 100.375 167.145 100.545 167.315 ;
        RECT 100.835 167.145 101.005 167.315 ;
        RECT 101.295 167.145 101.465 167.315 ;
        RECT 101.755 167.145 101.925 167.315 ;
        RECT 102.215 167.145 102.385 167.315 ;
        RECT 102.675 167.145 102.845 167.315 ;
        RECT 103.135 167.145 103.305 167.315 ;
        RECT 103.595 167.145 103.765 167.315 ;
        RECT 104.055 167.145 104.225 167.315 ;
        RECT 104.515 167.145 104.685 167.315 ;
        RECT 104.975 167.145 105.145 167.315 ;
        RECT 105.435 167.145 105.605 167.315 ;
        RECT 105.895 167.145 106.065 167.315 ;
        RECT 106.355 167.145 106.525 167.315 ;
        RECT 106.815 167.145 106.985 167.315 ;
        RECT 107.275 167.145 107.445 167.315 ;
        RECT 107.735 167.145 107.905 167.315 ;
        RECT 108.195 167.145 108.365 167.315 ;
        RECT 108.655 167.145 108.825 167.315 ;
        RECT 109.115 167.145 109.285 167.315 ;
        RECT 109.575 167.145 109.745 167.315 ;
        RECT 110.035 167.145 110.205 167.315 ;
        RECT 110.495 167.145 110.665 167.315 ;
        RECT 110.955 167.145 111.125 167.315 ;
        RECT 111.415 167.145 111.585 167.315 ;
        RECT 111.875 167.145 112.045 167.315 ;
        RECT 112.335 167.145 112.505 167.315 ;
        RECT 112.795 167.145 112.965 167.315 ;
        RECT 113.255 167.145 113.425 167.315 ;
        RECT 113.715 167.145 113.885 167.315 ;
        RECT 114.175 167.145 114.345 167.315 ;
        RECT 114.635 167.145 114.805 167.315 ;
        RECT 115.095 167.145 115.265 167.315 ;
        RECT 115.555 167.145 115.725 167.315 ;
        RECT 116.015 167.145 116.185 167.315 ;
        RECT 116.475 167.145 116.645 167.315 ;
        RECT 116.935 167.145 117.105 167.315 ;
        RECT 117.395 167.145 117.565 167.315 ;
        RECT 117.855 167.145 118.025 167.315 ;
        RECT 118.315 167.145 118.485 167.315 ;
        RECT 118.775 167.145 118.945 167.315 ;
        RECT 119.235 167.145 119.405 167.315 ;
        RECT 75.075 166.635 75.245 166.805 ;
        RECT 76.915 165.955 77.085 166.125 ;
        RECT 76.455 165.615 76.625 165.785 ;
        RECT 77.835 166.295 78.005 166.465 ;
        RECT 80.135 165.955 80.305 166.125 ;
        RECT 79.675 165.615 79.845 165.785 ;
        RECT 82.435 165.955 82.605 166.125 ;
        RECT 81.975 165.615 82.145 165.785 ;
        RECT 83.815 165.955 83.985 166.125 ;
        RECT 86.115 165.955 86.285 166.125 ;
        RECT 89.335 164.935 89.505 165.105 ;
        RECT 93.015 165.615 93.185 165.785 ;
        RECT 93.475 165.615 93.645 165.785 ;
        RECT 93.940 165.615 94.110 165.785 ;
        RECT 92.095 164.935 92.265 165.105 ;
        RECT 94.345 166.295 94.515 166.465 ;
        RECT 94.855 165.955 95.025 166.125 ;
        RECT 96.235 166.295 96.405 166.465 ;
        RECT 95.775 165.615 95.945 165.785 ;
        RECT 99.355 166.295 99.525 166.465 ;
        RECT 97.495 165.275 97.665 165.445 ;
        RECT 99.355 165.615 99.525 165.785 ;
        RECT 102.215 166.635 102.385 166.805 ;
        RECT 100.435 165.590 100.605 165.760 ;
        RECT 100.735 165.275 100.905 165.445 ;
        RECT 107.735 166.635 107.905 166.805 ;
        RECT 109.115 165.615 109.285 165.785 ;
        RECT 106.815 164.935 106.985 165.105 ;
        RECT 111.875 164.935 112.045 165.105 ;
        RECT 114.635 165.615 114.805 165.785 ;
        RECT 115.555 165.615 115.725 165.785 ;
        RECT 116.475 165.615 116.645 165.785 ;
        RECT 115.555 164.935 115.725 165.105 ;
        RECT 71.395 164.425 71.565 164.595 ;
        RECT 71.855 164.425 72.025 164.595 ;
        RECT 72.315 164.425 72.485 164.595 ;
        RECT 72.775 164.425 72.945 164.595 ;
        RECT 73.235 164.425 73.405 164.595 ;
        RECT 73.695 164.425 73.865 164.595 ;
        RECT 74.155 164.425 74.325 164.595 ;
        RECT 74.615 164.425 74.785 164.595 ;
        RECT 75.075 164.425 75.245 164.595 ;
        RECT 75.535 164.425 75.705 164.595 ;
        RECT 75.995 164.425 76.165 164.595 ;
        RECT 76.455 164.425 76.625 164.595 ;
        RECT 76.915 164.425 77.085 164.595 ;
        RECT 77.375 164.425 77.545 164.595 ;
        RECT 77.835 164.425 78.005 164.595 ;
        RECT 78.295 164.425 78.465 164.595 ;
        RECT 78.755 164.425 78.925 164.595 ;
        RECT 79.215 164.425 79.385 164.595 ;
        RECT 79.675 164.425 79.845 164.595 ;
        RECT 80.135 164.425 80.305 164.595 ;
        RECT 80.595 164.425 80.765 164.595 ;
        RECT 81.055 164.425 81.225 164.595 ;
        RECT 81.515 164.425 81.685 164.595 ;
        RECT 81.975 164.425 82.145 164.595 ;
        RECT 82.435 164.425 82.605 164.595 ;
        RECT 82.895 164.425 83.065 164.595 ;
        RECT 83.355 164.425 83.525 164.595 ;
        RECT 83.815 164.425 83.985 164.595 ;
        RECT 84.275 164.425 84.445 164.595 ;
        RECT 84.735 164.425 84.905 164.595 ;
        RECT 85.195 164.425 85.365 164.595 ;
        RECT 85.655 164.425 85.825 164.595 ;
        RECT 86.115 164.425 86.285 164.595 ;
        RECT 86.575 164.425 86.745 164.595 ;
        RECT 87.035 164.425 87.205 164.595 ;
        RECT 87.495 164.425 87.665 164.595 ;
        RECT 87.955 164.425 88.125 164.595 ;
        RECT 88.415 164.425 88.585 164.595 ;
        RECT 88.875 164.425 89.045 164.595 ;
        RECT 89.335 164.425 89.505 164.595 ;
        RECT 89.795 164.425 89.965 164.595 ;
        RECT 90.255 164.425 90.425 164.595 ;
        RECT 90.715 164.425 90.885 164.595 ;
        RECT 91.175 164.425 91.345 164.595 ;
        RECT 91.635 164.425 91.805 164.595 ;
        RECT 92.095 164.425 92.265 164.595 ;
        RECT 92.555 164.425 92.725 164.595 ;
        RECT 93.015 164.425 93.185 164.595 ;
        RECT 93.475 164.425 93.645 164.595 ;
        RECT 93.935 164.425 94.105 164.595 ;
        RECT 94.395 164.425 94.565 164.595 ;
        RECT 94.855 164.425 95.025 164.595 ;
        RECT 95.315 164.425 95.485 164.595 ;
        RECT 95.775 164.425 95.945 164.595 ;
        RECT 96.235 164.425 96.405 164.595 ;
        RECT 96.695 164.425 96.865 164.595 ;
        RECT 97.155 164.425 97.325 164.595 ;
        RECT 97.615 164.425 97.785 164.595 ;
        RECT 98.075 164.425 98.245 164.595 ;
        RECT 98.535 164.425 98.705 164.595 ;
        RECT 98.995 164.425 99.165 164.595 ;
        RECT 99.455 164.425 99.625 164.595 ;
        RECT 99.915 164.425 100.085 164.595 ;
        RECT 100.375 164.425 100.545 164.595 ;
        RECT 100.835 164.425 101.005 164.595 ;
        RECT 101.295 164.425 101.465 164.595 ;
        RECT 101.755 164.425 101.925 164.595 ;
        RECT 102.215 164.425 102.385 164.595 ;
        RECT 102.675 164.425 102.845 164.595 ;
        RECT 103.135 164.425 103.305 164.595 ;
        RECT 103.595 164.425 103.765 164.595 ;
        RECT 104.055 164.425 104.225 164.595 ;
        RECT 104.515 164.425 104.685 164.595 ;
        RECT 104.975 164.425 105.145 164.595 ;
        RECT 105.435 164.425 105.605 164.595 ;
        RECT 105.895 164.425 106.065 164.595 ;
        RECT 106.355 164.425 106.525 164.595 ;
        RECT 106.815 164.425 106.985 164.595 ;
        RECT 107.275 164.425 107.445 164.595 ;
        RECT 107.735 164.425 107.905 164.595 ;
        RECT 108.195 164.425 108.365 164.595 ;
        RECT 108.655 164.425 108.825 164.595 ;
        RECT 109.115 164.425 109.285 164.595 ;
        RECT 109.575 164.425 109.745 164.595 ;
        RECT 110.035 164.425 110.205 164.595 ;
        RECT 110.495 164.425 110.665 164.595 ;
        RECT 110.955 164.425 111.125 164.595 ;
        RECT 111.415 164.425 111.585 164.595 ;
        RECT 111.875 164.425 112.045 164.595 ;
        RECT 112.335 164.425 112.505 164.595 ;
        RECT 112.795 164.425 112.965 164.595 ;
        RECT 113.255 164.425 113.425 164.595 ;
        RECT 113.715 164.425 113.885 164.595 ;
        RECT 114.175 164.425 114.345 164.595 ;
        RECT 114.635 164.425 114.805 164.595 ;
        RECT 115.095 164.425 115.265 164.595 ;
        RECT 115.555 164.425 115.725 164.595 ;
        RECT 116.015 164.425 116.185 164.595 ;
        RECT 116.475 164.425 116.645 164.595 ;
        RECT 116.935 164.425 117.105 164.595 ;
        RECT 117.395 164.425 117.565 164.595 ;
        RECT 117.855 164.425 118.025 164.595 ;
        RECT 118.315 164.425 118.485 164.595 ;
        RECT 118.775 164.425 118.945 164.595 ;
        RECT 119.235 164.425 119.405 164.595 ;
        RECT 75.535 162.895 75.705 163.065 ;
        RECT 76.000 163.235 76.170 163.405 ;
        RECT 76.915 162.895 77.085 163.065 ;
        RECT 76.405 162.555 76.575 162.725 ;
        RECT 77.835 163.235 78.005 163.405 ;
        RECT 79.195 163.575 79.365 163.745 ;
        RECT 79.555 163.575 79.725 163.745 ;
        RECT 78.295 162.555 78.465 162.725 ;
        RECT 81.415 163.235 81.585 163.405 ;
        RECT 82.795 163.575 82.965 163.745 ;
        RECT 82.495 163.260 82.665 163.430 ;
        RECT 81.415 162.555 81.585 162.725 ;
        RECT 84.275 162.215 84.445 162.385 ;
        RECT 85.655 163.915 85.825 164.085 ;
        RECT 87.135 163.575 87.305 163.745 ;
        RECT 87.435 163.260 87.605 163.430 ;
        RECT 88.515 163.235 88.685 163.405 ;
        RECT 90.375 163.575 90.545 163.745 ;
        RECT 90.735 163.575 90.905 163.745 ;
        RECT 88.515 162.555 88.685 162.725 ;
        RECT 92.095 163.235 92.265 163.405 ;
        RECT 91.635 162.555 91.805 162.725 ;
        RECT 93.015 163.575 93.185 163.745 ;
        RECT 93.525 162.555 93.695 162.725 ;
        RECT 93.930 163.235 94.100 163.405 ;
        RECT 94.395 162.895 94.565 163.065 ;
        RECT 97.615 162.895 97.785 163.065 ;
        RECT 98.080 163.235 98.250 163.405 ;
        RECT 98.995 163.575 99.165 163.745 ;
        RECT 98.485 162.555 98.655 162.725 ;
        RECT 99.915 163.235 100.085 163.405 ;
        RECT 101.275 163.575 101.445 163.745 ;
        RECT 101.635 163.575 101.805 163.745 ;
        RECT 100.375 162.555 100.545 162.725 ;
        RECT 103.495 163.235 103.665 163.405 ;
        RECT 104.875 163.575 105.045 163.745 ;
        RECT 104.575 163.260 104.745 163.430 ;
        RECT 103.495 162.555 103.665 162.725 ;
        RECT 106.355 162.215 106.525 162.385 ;
        RECT 108.195 162.895 108.365 163.065 ;
        RECT 108.680 162.555 108.850 162.725 ;
        RECT 109.075 162.895 109.245 163.065 ;
        RECT 109.530 163.575 109.700 163.745 ;
        RECT 110.265 162.895 110.435 163.065 ;
        RECT 110.780 162.555 110.950 162.725 ;
        RECT 112.350 162.555 112.520 162.725 ;
        RECT 112.785 162.895 112.955 163.065 ;
        RECT 115.095 162.215 115.265 162.385 ;
        RECT 71.395 161.705 71.565 161.875 ;
        RECT 71.855 161.705 72.025 161.875 ;
        RECT 72.315 161.705 72.485 161.875 ;
        RECT 72.775 161.705 72.945 161.875 ;
        RECT 73.235 161.705 73.405 161.875 ;
        RECT 73.695 161.705 73.865 161.875 ;
        RECT 74.155 161.705 74.325 161.875 ;
        RECT 74.615 161.705 74.785 161.875 ;
        RECT 75.075 161.705 75.245 161.875 ;
        RECT 75.535 161.705 75.705 161.875 ;
        RECT 75.995 161.705 76.165 161.875 ;
        RECT 76.455 161.705 76.625 161.875 ;
        RECT 76.915 161.705 77.085 161.875 ;
        RECT 77.375 161.705 77.545 161.875 ;
        RECT 77.835 161.705 78.005 161.875 ;
        RECT 78.295 161.705 78.465 161.875 ;
        RECT 78.755 161.705 78.925 161.875 ;
        RECT 79.215 161.705 79.385 161.875 ;
        RECT 79.675 161.705 79.845 161.875 ;
        RECT 80.135 161.705 80.305 161.875 ;
        RECT 80.595 161.705 80.765 161.875 ;
        RECT 81.055 161.705 81.225 161.875 ;
        RECT 81.515 161.705 81.685 161.875 ;
        RECT 81.975 161.705 82.145 161.875 ;
        RECT 82.435 161.705 82.605 161.875 ;
        RECT 82.895 161.705 83.065 161.875 ;
        RECT 83.355 161.705 83.525 161.875 ;
        RECT 83.815 161.705 83.985 161.875 ;
        RECT 84.275 161.705 84.445 161.875 ;
        RECT 84.735 161.705 84.905 161.875 ;
        RECT 85.195 161.705 85.365 161.875 ;
        RECT 85.655 161.705 85.825 161.875 ;
        RECT 86.115 161.705 86.285 161.875 ;
        RECT 86.575 161.705 86.745 161.875 ;
        RECT 87.035 161.705 87.205 161.875 ;
        RECT 87.495 161.705 87.665 161.875 ;
        RECT 87.955 161.705 88.125 161.875 ;
        RECT 88.415 161.705 88.585 161.875 ;
        RECT 88.875 161.705 89.045 161.875 ;
        RECT 89.335 161.705 89.505 161.875 ;
        RECT 89.795 161.705 89.965 161.875 ;
        RECT 90.255 161.705 90.425 161.875 ;
        RECT 90.715 161.705 90.885 161.875 ;
        RECT 91.175 161.705 91.345 161.875 ;
        RECT 91.635 161.705 91.805 161.875 ;
        RECT 92.095 161.705 92.265 161.875 ;
        RECT 92.555 161.705 92.725 161.875 ;
        RECT 93.015 161.705 93.185 161.875 ;
        RECT 93.475 161.705 93.645 161.875 ;
        RECT 93.935 161.705 94.105 161.875 ;
        RECT 94.395 161.705 94.565 161.875 ;
        RECT 94.855 161.705 95.025 161.875 ;
        RECT 95.315 161.705 95.485 161.875 ;
        RECT 95.775 161.705 95.945 161.875 ;
        RECT 96.235 161.705 96.405 161.875 ;
        RECT 96.695 161.705 96.865 161.875 ;
        RECT 97.155 161.705 97.325 161.875 ;
        RECT 97.615 161.705 97.785 161.875 ;
        RECT 98.075 161.705 98.245 161.875 ;
        RECT 98.535 161.705 98.705 161.875 ;
        RECT 98.995 161.705 99.165 161.875 ;
        RECT 99.455 161.705 99.625 161.875 ;
        RECT 99.915 161.705 100.085 161.875 ;
        RECT 100.375 161.705 100.545 161.875 ;
        RECT 100.835 161.705 101.005 161.875 ;
        RECT 101.295 161.705 101.465 161.875 ;
        RECT 101.755 161.705 101.925 161.875 ;
        RECT 102.215 161.705 102.385 161.875 ;
        RECT 102.675 161.705 102.845 161.875 ;
        RECT 103.135 161.705 103.305 161.875 ;
        RECT 103.595 161.705 103.765 161.875 ;
        RECT 104.055 161.705 104.225 161.875 ;
        RECT 104.515 161.705 104.685 161.875 ;
        RECT 104.975 161.705 105.145 161.875 ;
        RECT 105.435 161.705 105.605 161.875 ;
        RECT 105.895 161.705 106.065 161.875 ;
        RECT 106.355 161.705 106.525 161.875 ;
        RECT 106.815 161.705 106.985 161.875 ;
        RECT 107.275 161.705 107.445 161.875 ;
        RECT 107.735 161.705 107.905 161.875 ;
        RECT 108.195 161.705 108.365 161.875 ;
        RECT 108.655 161.705 108.825 161.875 ;
        RECT 109.115 161.705 109.285 161.875 ;
        RECT 109.575 161.705 109.745 161.875 ;
        RECT 110.035 161.705 110.205 161.875 ;
        RECT 110.495 161.705 110.665 161.875 ;
        RECT 110.955 161.705 111.125 161.875 ;
        RECT 111.415 161.705 111.585 161.875 ;
        RECT 111.875 161.705 112.045 161.875 ;
        RECT 112.335 161.705 112.505 161.875 ;
        RECT 112.795 161.705 112.965 161.875 ;
        RECT 113.255 161.705 113.425 161.875 ;
        RECT 113.715 161.705 113.885 161.875 ;
        RECT 114.175 161.705 114.345 161.875 ;
        RECT 114.635 161.705 114.805 161.875 ;
        RECT 115.095 161.705 115.265 161.875 ;
        RECT 115.555 161.705 115.725 161.875 ;
        RECT 116.015 161.705 116.185 161.875 ;
        RECT 116.475 161.705 116.645 161.875 ;
        RECT 116.935 161.705 117.105 161.875 ;
        RECT 117.395 161.705 117.565 161.875 ;
        RECT 117.855 161.705 118.025 161.875 ;
        RECT 118.315 161.705 118.485 161.875 ;
        RECT 118.775 161.705 118.945 161.875 ;
        RECT 119.235 161.705 119.405 161.875 ;
        RECT 86.575 160.515 86.745 160.685 ;
        RECT 87.955 160.175 88.125 160.345 ;
        RECT 102.215 160.175 102.385 160.345 ;
        RECT 105.435 159.495 105.605 159.665 ;
        RECT 105.895 160.175 106.065 160.345 ;
        RECT 111.415 160.515 111.585 160.685 ;
        RECT 108.655 160.175 108.825 160.345 ;
        RECT 110.495 160.175 110.665 160.345 ;
        RECT 111.875 161.195 112.045 161.365 ;
        RECT 112.335 160.855 112.505 161.025 ;
        RECT 114.175 161.195 114.345 161.365 ;
        RECT 112.795 160.175 112.965 160.345 ;
        RECT 114.635 160.175 114.805 160.345 ;
        RECT 117.395 160.515 117.565 160.685 ;
        RECT 71.395 158.985 71.565 159.155 ;
        RECT 71.855 158.985 72.025 159.155 ;
        RECT 72.315 158.985 72.485 159.155 ;
        RECT 72.775 158.985 72.945 159.155 ;
        RECT 73.235 158.985 73.405 159.155 ;
        RECT 73.695 158.985 73.865 159.155 ;
        RECT 74.155 158.985 74.325 159.155 ;
        RECT 74.615 158.985 74.785 159.155 ;
        RECT 75.075 158.985 75.245 159.155 ;
        RECT 75.535 158.985 75.705 159.155 ;
        RECT 75.995 158.985 76.165 159.155 ;
        RECT 76.455 158.985 76.625 159.155 ;
        RECT 76.915 158.985 77.085 159.155 ;
        RECT 77.375 158.985 77.545 159.155 ;
        RECT 77.835 158.985 78.005 159.155 ;
        RECT 78.295 158.985 78.465 159.155 ;
        RECT 78.755 158.985 78.925 159.155 ;
        RECT 79.215 158.985 79.385 159.155 ;
        RECT 79.675 158.985 79.845 159.155 ;
        RECT 80.135 158.985 80.305 159.155 ;
        RECT 80.595 158.985 80.765 159.155 ;
        RECT 81.055 158.985 81.225 159.155 ;
        RECT 81.515 158.985 81.685 159.155 ;
        RECT 81.975 158.985 82.145 159.155 ;
        RECT 82.435 158.985 82.605 159.155 ;
        RECT 82.895 158.985 83.065 159.155 ;
        RECT 83.355 158.985 83.525 159.155 ;
        RECT 83.815 158.985 83.985 159.155 ;
        RECT 84.275 158.985 84.445 159.155 ;
        RECT 84.735 158.985 84.905 159.155 ;
        RECT 85.195 158.985 85.365 159.155 ;
        RECT 85.655 158.985 85.825 159.155 ;
        RECT 86.115 158.985 86.285 159.155 ;
        RECT 86.575 158.985 86.745 159.155 ;
        RECT 87.035 158.985 87.205 159.155 ;
        RECT 87.495 158.985 87.665 159.155 ;
        RECT 87.955 158.985 88.125 159.155 ;
        RECT 88.415 158.985 88.585 159.155 ;
        RECT 88.875 158.985 89.045 159.155 ;
        RECT 89.335 158.985 89.505 159.155 ;
        RECT 89.795 158.985 89.965 159.155 ;
        RECT 90.255 158.985 90.425 159.155 ;
        RECT 90.715 158.985 90.885 159.155 ;
        RECT 91.175 158.985 91.345 159.155 ;
        RECT 91.635 158.985 91.805 159.155 ;
        RECT 92.095 158.985 92.265 159.155 ;
        RECT 92.555 158.985 92.725 159.155 ;
        RECT 93.015 158.985 93.185 159.155 ;
        RECT 93.475 158.985 93.645 159.155 ;
        RECT 93.935 158.985 94.105 159.155 ;
        RECT 94.395 158.985 94.565 159.155 ;
        RECT 94.855 158.985 95.025 159.155 ;
        RECT 95.315 158.985 95.485 159.155 ;
        RECT 95.775 158.985 95.945 159.155 ;
        RECT 96.235 158.985 96.405 159.155 ;
        RECT 96.695 158.985 96.865 159.155 ;
        RECT 97.155 158.985 97.325 159.155 ;
        RECT 97.615 158.985 97.785 159.155 ;
        RECT 98.075 158.985 98.245 159.155 ;
        RECT 98.535 158.985 98.705 159.155 ;
        RECT 98.995 158.985 99.165 159.155 ;
        RECT 99.455 158.985 99.625 159.155 ;
        RECT 99.915 158.985 100.085 159.155 ;
        RECT 100.375 158.985 100.545 159.155 ;
        RECT 100.835 158.985 101.005 159.155 ;
        RECT 101.295 158.985 101.465 159.155 ;
        RECT 101.755 158.985 101.925 159.155 ;
        RECT 102.215 158.985 102.385 159.155 ;
        RECT 102.675 158.985 102.845 159.155 ;
        RECT 103.135 158.985 103.305 159.155 ;
        RECT 103.595 158.985 103.765 159.155 ;
        RECT 104.055 158.985 104.225 159.155 ;
        RECT 104.515 158.985 104.685 159.155 ;
        RECT 104.975 158.985 105.145 159.155 ;
        RECT 105.435 158.985 105.605 159.155 ;
        RECT 105.895 158.985 106.065 159.155 ;
        RECT 106.355 158.985 106.525 159.155 ;
        RECT 106.815 158.985 106.985 159.155 ;
        RECT 107.275 158.985 107.445 159.155 ;
        RECT 107.735 158.985 107.905 159.155 ;
        RECT 108.195 158.985 108.365 159.155 ;
        RECT 108.655 158.985 108.825 159.155 ;
        RECT 109.115 158.985 109.285 159.155 ;
        RECT 109.575 158.985 109.745 159.155 ;
        RECT 110.035 158.985 110.205 159.155 ;
        RECT 110.495 158.985 110.665 159.155 ;
        RECT 110.955 158.985 111.125 159.155 ;
        RECT 111.415 158.985 111.585 159.155 ;
        RECT 111.875 158.985 112.045 159.155 ;
        RECT 112.335 158.985 112.505 159.155 ;
        RECT 112.795 158.985 112.965 159.155 ;
        RECT 113.255 158.985 113.425 159.155 ;
        RECT 113.715 158.985 113.885 159.155 ;
        RECT 114.175 158.985 114.345 159.155 ;
        RECT 114.635 158.985 114.805 159.155 ;
        RECT 115.095 158.985 115.265 159.155 ;
        RECT 115.555 158.985 115.725 159.155 ;
        RECT 116.015 158.985 116.185 159.155 ;
        RECT 116.475 158.985 116.645 159.155 ;
        RECT 116.935 158.985 117.105 159.155 ;
        RECT 117.395 158.985 117.565 159.155 ;
        RECT 117.855 158.985 118.025 159.155 ;
        RECT 118.315 158.985 118.485 159.155 ;
        RECT 118.775 158.985 118.945 159.155 ;
        RECT 119.235 158.985 119.405 159.155 ;
        RECT 82.435 157.795 82.605 157.965 ;
        RECT 82.895 157.455 83.065 157.625 ;
        RECT 84.275 157.455 84.445 157.625 ;
        RECT 86.575 157.795 86.745 157.965 ;
        RECT 86.115 157.455 86.285 157.625 ;
        RECT 84.735 156.775 84.905 156.945 ;
        RECT 88.875 157.795 89.045 157.965 ;
        RECT 88.415 157.455 88.585 157.625 ;
        RECT 90.715 157.455 90.885 157.625 ;
        RECT 91.635 157.455 91.805 157.625 ;
        RECT 101.755 158.475 101.925 158.645 ;
        RECT 94.855 156.775 95.025 156.945 ;
        RECT 106.355 158.475 106.525 158.645 ;
        RECT 103.135 157.795 103.305 157.965 ;
        RECT 103.595 157.795 103.765 157.965 ;
        RECT 104.055 157.455 104.225 157.625 ;
        RECT 105.435 157.795 105.605 157.965 ;
        RECT 104.515 156.775 104.685 156.945 ;
        RECT 107.730 158.135 107.900 158.305 ;
        RECT 108.145 157.115 108.315 157.285 ;
        RECT 109.575 157.795 109.745 157.965 ;
        RECT 110.955 157.455 111.125 157.625 ;
        RECT 113.250 157.795 113.420 157.965 ;
        RECT 111.375 157.115 111.545 157.285 ;
        RECT 112.335 157.115 112.505 157.285 ;
        RECT 114.635 157.795 114.805 157.965 ;
        RECT 115.555 157.455 115.725 157.625 ;
        RECT 71.395 156.265 71.565 156.435 ;
        RECT 71.855 156.265 72.025 156.435 ;
        RECT 72.315 156.265 72.485 156.435 ;
        RECT 72.775 156.265 72.945 156.435 ;
        RECT 73.235 156.265 73.405 156.435 ;
        RECT 73.695 156.265 73.865 156.435 ;
        RECT 74.155 156.265 74.325 156.435 ;
        RECT 74.615 156.265 74.785 156.435 ;
        RECT 75.075 156.265 75.245 156.435 ;
        RECT 75.535 156.265 75.705 156.435 ;
        RECT 75.995 156.265 76.165 156.435 ;
        RECT 76.455 156.265 76.625 156.435 ;
        RECT 76.915 156.265 77.085 156.435 ;
        RECT 77.375 156.265 77.545 156.435 ;
        RECT 77.835 156.265 78.005 156.435 ;
        RECT 78.295 156.265 78.465 156.435 ;
        RECT 78.755 156.265 78.925 156.435 ;
        RECT 79.215 156.265 79.385 156.435 ;
        RECT 79.675 156.265 79.845 156.435 ;
        RECT 80.135 156.265 80.305 156.435 ;
        RECT 80.595 156.265 80.765 156.435 ;
        RECT 81.055 156.265 81.225 156.435 ;
        RECT 81.515 156.265 81.685 156.435 ;
        RECT 81.975 156.265 82.145 156.435 ;
        RECT 82.435 156.265 82.605 156.435 ;
        RECT 82.895 156.265 83.065 156.435 ;
        RECT 83.355 156.265 83.525 156.435 ;
        RECT 83.815 156.265 83.985 156.435 ;
        RECT 84.275 156.265 84.445 156.435 ;
        RECT 84.735 156.265 84.905 156.435 ;
        RECT 85.195 156.265 85.365 156.435 ;
        RECT 85.655 156.265 85.825 156.435 ;
        RECT 86.115 156.265 86.285 156.435 ;
        RECT 86.575 156.265 86.745 156.435 ;
        RECT 87.035 156.265 87.205 156.435 ;
        RECT 87.495 156.265 87.665 156.435 ;
        RECT 87.955 156.265 88.125 156.435 ;
        RECT 88.415 156.265 88.585 156.435 ;
        RECT 88.875 156.265 89.045 156.435 ;
        RECT 89.335 156.265 89.505 156.435 ;
        RECT 89.795 156.265 89.965 156.435 ;
        RECT 90.255 156.265 90.425 156.435 ;
        RECT 90.715 156.265 90.885 156.435 ;
        RECT 91.175 156.265 91.345 156.435 ;
        RECT 91.635 156.265 91.805 156.435 ;
        RECT 92.095 156.265 92.265 156.435 ;
        RECT 92.555 156.265 92.725 156.435 ;
        RECT 93.015 156.265 93.185 156.435 ;
        RECT 93.475 156.265 93.645 156.435 ;
        RECT 93.935 156.265 94.105 156.435 ;
        RECT 94.395 156.265 94.565 156.435 ;
        RECT 94.855 156.265 95.025 156.435 ;
        RECT 95.315 156.265 95.485 156.435 ;
        RECT 95.775 156.265 95.945 156.435 ;
        RECT 96.235 156.265 96.405 156.435 ;
        RECT 96.695 156.265 96.865 156.435 ;
        RECT 97.155 156.265 97.325 156.435 ;
        RECT 97.615 156.265 97.785 156.435 ;
        RECT 98.075 156.265 98.245 156.435 ;
        RECT 98.535 156.265 98.705 156.435 ;
        RECT 98.995 156.265 99.165 156.435 ;
        RECT 99.455 156.265 99.625 156.435 ;
        RECT 99.915 156.265 100.085 156.435 ;
        RECT 100.375 156.265 100.545 156.435 ;
        RECT 100.835 156.265 101.005 156.435 ;
        RECT 101.295 156.265 101.465 156.435 ;
        RECT 101.755 156.265 101.925 156.435 ;
        RECT 102.215 156.265 102.385 156.435 ;
        RECT 102.675 156.265 102.845 156.435 ;
        RECT 103.135 156.265 103.305 156.435 ;
        RECT 103.595 156.265 103.765 156.435 ;
        RECT 104.055 156.265 104.225 156.435 ;
        RECT 104.515 156.265 104.685 156.435 ;
        RECT 104.975 156.265 105.145 156.435 ;
        RECT 105.435 156.265 105.605 156.435 ;
        RECT 105.895 156.265 106.065 156.435 ;
        RECT 106.355 156.265 106.525 156.435 ;
        RECT 106.815 156.265 106.985 156.435 ;
        RECT 107.275 156.265 107.445 156.435 ;
        RECT 107.735 156.265 107.905 156.435 ;
        RECT 108.195 156.265 108.365 156.435 ;
        RECT 108.655 156.265 108.825 156.435 ;
        RECT 109.115 156.265 109.285 156.435 ;
        RECT 109.575 156.265 109.745 156.435 ;
        RECT 110.035 156.265 110.205 156.435 ;
        RECT 110.495 156.265 110.665 156.435 ;
        RECT 110.955 156.265 111.125 156.435 ;
        RECT 111.415 156.265 111.585 156.435 ;
        RECT 111.875 156.265 112.045 156.435 ;
        RECT 112.335 156.265 112.505 156.435 ;
        RECT 112.795 156.265 112.965 156.435 ;
        RECT 113.255 156.265 113.425 156.435 ;
        RECT 113.715 156.265 113.885 156.435 ;
        RECT 114.175 156.265 114.345 156.435 ;
        RECT 114.635 156.265 114.805 156.435 ;
        RECT 115.095 156.265 115.265 156.435 ;
        RECT 115.555 156.265 115.725 156.435 ;
        RECT 116.015 156.265 116.185 156.435 ;
        RECT 116.475 156.265 116.645 156.435 ;
        RECT 116.935 156.265 117.105 156.435 ;
        RECT 117.395 156.265 117.565 156.435 ;
        RECT 117.855 156.265 118.025 156.435 ;
        RECT 118.315 156.265 118.485 156.435 ;
        RECT 118.775 156.265 118.945 156.435 ;
        RECT 119.235 156.265 119.405 156.435 ;
        RECT 73.695 155.075 73.865 155.245 ;
        RECT 74.160 154.735 74.330 154.905 ;
        RECT 74.565 155.415 74.735 155.585 ;
        RECT 75.075 154.395 75.245 154.565 ;
        RECT 76.455 155.415 76.625 155.585 ;
        RECT 75.995 154.735 76.165 154.905 ;
        RECT 79.575 155.415 79.745 155.585 ;
        RECT 77.715 154.395 77.885 154.565 ;
        RECT 79.575 154.735 79.745 154.905 ;
        RECT 80.655 154.710 80.825 154.880 ;
        RECT 80.955 154.395 81.125 154.565 ;
        RECT 82.435 154.055 82.605 154.225 ;
        RECT 84.735 154.055 84.905 154.225 ;
        RECT 88.415 155.755 88.585 155.925 ;
        RECT 87.495 154.735 87.665 154.905 ;
        RECT 91.635 154.735 91.805 154.905 ;
        RECT 92.095 155.075 92.265 155.245 ;
        RECT 92.560 154.735 92.730 154.905 ;
        RECT 92.965 155.415 93.135 155.585 ;
        RECT 93.410 155.755 93.580 155.925 ;
        RECT 94.855 155.415 95.025 155.585 ;
        RECT 94.395 154.735 94.565 154.905 ;
        RECT 97.975 155.415 98.145 155.585 ;
        RECT 96.115 154.395 96.285 154.565 ;
        RECT 97.975 154.735 98.145 154.905 ;
        RECT 100.835 155.755 101.005 155.925 ;
        RECT 101.780 155.415 101.950 155.585 ;
        RECT 99.055 154.710 99.225 154.880 ;
        RECT 99.355 154.395 99.525 154.565 ;
        RECT 101.295 155.075 101.465 155.245 ;
        RECT 102.175 155.075 102.345 155.245 ;
        RECT 102.630 154.395 102.800 154.565 ;
        RECT 103.880 155.415 104.050 155.585 ;
        RECT 103.365 155.075 103.535 155.245 ;
        RECT 105.450 155.415 105.620 155.585 ;
        RECT 105.885 155.075 106.055 155.245 ;
        RECT 108.195 155.755 108.365 155.925 ;
        RECT 109.115 155.415 109.285 155.585 ;
        RECT 111.440 155.415 111.610 155.585 ;
        RECT 110.955 155.075 111.125 155.245 ;
        RECT 109.575 154.735 109.745 154.905 ;
        RECT 111.835 155.075 112.005 155.245 ;
        RECT 112.290 154.395 112.460 154.565 ;
        RECT 113.540 155.415 113.710 155.585 ;
        RECT 113.025 155.075 113.195 155.245 ;
        RECT 115.110 155.415 115.280 155.585 ;
        RECT 115.545 155.075 115.715 155.245 ;
        RECT 117.855 155.755 118.025 155.925 ;
        RECT 71.395 153.545 71.565 153.715 ;
        RECT 71.855 153.545 72.025 153.715 ;
        RECT 72.315 153.545 72.485 153.715 ;
        RECT 72.775 153.545 72.945 153.715 ;
        RECT 73.235 153.545 73.405 153.715 ;
        RECT 73.695 153.545 73.865 153.715 ;
        RECT 74.155 153.545 74.325 153.715 ;
        RECT 74.615 153.545 74.785 153.715 ;
        RECT 75.075 153.545 75.245 153.715 ;
        RECT 75.535 153.545 75.705 153.715 ;
        RECT 75.995 153.545 76.165 153.715 ;
        RECT 76.455 153.545 76.625 153.715 ;
        RECT 76.915 153.545 77.085 153.715 ;
        RECT 77.375 153.545 77.545 153.715 ;
        RECT 77.835 153.545 78.005 153.715 ;
        RECT 78.295 153.545 78.465 153.715 ;
        RECT 78.755 153.545 78.925 153.715 ;
        RECT 79.215 153.545 79.385 153.715 ;
        RECT 79.675 153.545 79.845 153.715 ;
        RECT 80.135 153.545 80.305 153.715 ;
        RECT 80.595 153.545 80.765 153.715 ;
        RECT 81.055 153.545 81.225 153.715 ;
        RECT 81.515 153.545 81.685 153.715 ;
        RECT 81.975 153.545 82.145 153.715 ;
        RECT 82.435 153.545 82.605 153.715 ;
        RECT 82.895 153.545 83.065 153.715 ;
        RECT 83.355 153.545 83.525 153.715 ;
        RECT 83.815 153.545 83.985 153.715 ;
        RECT 84.275 153.545 84.445 153.715 ;
        RECT 84.735 153.545 84.905 153.715 ;
        RECT 85.195 153.545 85.365 153.715 ;
        RECT 85.655 153.545 85.825 153.715 ;
        RECT 86.115 153.545 86.285 153.715 ;
        RECT 86.575 153.545 86.745 153.715 ;
        RECT 87.035 153.545 87.205 153.715 ;
        RECT 87.495 153.545 87.665 153.715 ;
        RECT 87.955 153.545 88.125 153.715 ;
        RECT 88.415 153.545 88.585 153.715 ;
        RECT 88.875 153.545 89.045 153.715 ;
        RECT 89.335 153.545 89.505 153.715 ;
        RECT 89.795 153.545 89.965 153.715 ;
        RECT 90.255 153.545 90.425 153.715 ;
        RECT 90.715 153.545 90.885 153.715 ;
        RECT 91.175 153.545 91.345 153.715 ;
        RECT 91.635 153.545 91.805 153.715 ;
        RECT 92.095 153.545 92.265 153.715 ;
        RECT 92.555 153.545 92.725 153.715 ;
        RECT 93.015 153.545 93.185 153.715 ;
        RECT 93.475 153.545 93.645 153.715 ;
        RECT 93.935 153.545 94.105 153.715 ;
        RECT 94.395 153.545 94.565 153.715 ;
        RECT 94.855 153.545 95.025 153.715 ;
        RECT 95.315 153.545 95.485 153.715 ;
        RECT 95.775 153.545 95.945 153.715 ;
        RECT 96.235 153.545 96.405 153.715 ;
        RECT 96.695 153.545 96.865 153.715 ;
        RECT 97.155 153.545 97.325 153.715 ;
        RECT 97.615 153.545 97.785 153.715 ;
        RECT 98.075 153.545 98.245 153.715 ;
        RECT 98.535 153.545 98.705 153.715 ;
        RECT 98.995 153.545 99.165 153.715 ;
        RECT 99.455 153.545 99.625 153.715 ;
        RECT 99.915 153.545 100.085 153.715 ;
        RECT 100.375 153.545 100.545 153.715 ;
        RECT 100.835 153.545 101.005 153.715 ;
        RECT 101.295 153.545 101.465 153.715 ;
        RECT 101.755 153.545 101.925 153.715 ;
        RECT 102.215 153.545 102.385 153.715 ;
        RECT 102.675 153.545 102.845 153.715 ;
        RECT 103.135 153.545 103.305 153.715 ;
        RECT 103.595 153.545 103.765 153.715 ;
        RECT 104.055 153.545 104.225 153.715 ;
        RECT 104.515 153.545 104.685 153.715 ;
        RECT 104.975 153.545 105.145 153.715 ;
        RECT 105.435 153.545 105.605 153.715 ;
        RECT 105.895 153.545 106.065 153.715 ;
        RECT 106.355 153.545 106.525 153.715 ;
        RECT 106.815 153.545 106.985 153.715 ;
        RECT 107.275 153.545 107.445 153.715 ;
        RECT 107.735 153.545 107.905 153.715 ;
        RECT 108.195 153.545 108.365 153.715 ;
        RECT 108.655 153.545 108.825 153.715 ;
        RECT 109.115 153.545 109.285 153.715 ;
        RECT 109.575 153.545 109.745 153.715 ;
        RECT 110.035 153.545 110.205 153.715 ;
        RECT 110.495 153.545 110.665 153.715 ;
        RECT 110.955 153.545 111.125 153.715 ;
        RECT 111.415 153.545 111.585 153.715 ;
        RECT 111.875 153.545 112.045 153.715 ;
        RECT 112.335 153.545 112.505 153.715 ;
        RECT 112.795 153.545 112.965 153.715 ;
        RECT 113.255 153.545 113.425 153.715 ;
        RECT 113.715 153.545 113.885 153.715 ;
        RECT 114.175 153.545 114.345 153.715 ;
        RECT 114.635 153.545 114.805 153.715 ;
        RECT 115.095 153.545 115.265 153.715 ;
        RECT 115.555 153.545 115.725 153.715 ;
        RECT 116.015 153.545 116.185 153.715 ;
        RECT 116.475 153.545 116.645 153.715 ;
        RECT 116.935 153.545 117.105 153.715 ;
        RECT 117.395 153.545 117.565 153.715 ;
        RECT 117.855 153.545 118.025 153.715 ;
        RECT 118.315 153.545 118.485 153.715 ;
        RECT 118.775 153.545 118.945 153.715 ;
        RECT 119.235 153.545 119.405 153.715 ;
        RECT 17.715 153.005 17.890 153.190 ;
        RECT 20.720 153.025 20.890 153.200 ;
        RECT 15.245 147.590 15.980 148.210 ;
        RECT 18.960 151.225 19.130 152.105 ;
        RECT 19.400 151.225 19.570 152.105 ;
        RECT 19.840 151.225 20.010 152.105 ;
        RECT 20.470 151.225 20.640 152.105 ;
        RECT 77.835 153.035 78.005 153.205 ;
        RECT 20.910 151.225 21.080 152.105 ;
        RECT 21.350 151.225 21.520 152.105 ;
        RECT 81.515 152.015 81.685 152.185 ;
        RECT 83.355 152.355 83.525 152.525 ;
        RECT 83.815 152.015 83.985 152.185 ;
        RECT 96.695 152.695 96.865 152.865 ;
        RECT 89.335 151.335 89.505 151.505 ;
        RECT 103.595 152.695 103.765 152.865 ;
        RECT 101.295 152.355 101.465 152.525 ;
        RECT 101.755 152.355 101.925 152.525 ;
        RECT 102.675 152.355 102.845 152.525 ;
        RECT 102.215 151.675 102.385 151.845 ;
        RECT 104.055 152.015 104.225 152.185 ;
        RECT 104.540 151.675 104.710 151.845 ;
        RECT 104.935 152.015 105.105 152.185 ;
        RECT 105.390 152.355 105.560 152.525 ;
        RECT 106.125 152.015 106.295 152.185 ;
        RECT 106.640 151.675 106.810 151.845 ;
        RECT 108.210 151.675 108.380 151.845 ;
        RECT 108.645 152.015 108.815 152.185 ;
        RECT 110.955 153.035 111.125 153.205 ;
        RECT 111.875 152.355 112.045 152.525 ;
        RECT 115.095 153.035 115.265 153.205 ;
        RECT 116.935 153.035 117.105 153.205 ;
        RECT 117.855 152.355 118.025 152.525 ;
        RECT 71.395 150.825 71.565 150.995 ;
        RECT 71.855 150.825 72.025 150.995 ;
        RECT 72.315 150.825 72.485 150.995 ;
        RECT 72.775 150.825 72.945 150.995 ;
        RECT 73.235 150.825 73.405 150.995 ;
        RECT 73.695 150.825 73.865 150.995 ;
        RECT 74.155 150.825 74.325 150.995 ;
        RECT 74.615 150.825 74.785 150.995 ;
        RECT 75.075 150.825 75.245 150.995 ;
        RECT 75.535 150.825 75.705 150.995 ;
        RECT 75.995 150.825 76.165 150.995 ;
        RECT 76.455 150.825 76.625 150.995 ;
        RECT 76.915 150.825 77.085 150.995 ;
        RECT 77.375 150.825 77.545 150.995 ;
        RECT 77.835 150.825 78.005 150.995 ;
        RECT 78.295 150.825 78.465 150.995 ;
        RECT 78.755 150.825 78.925 150.995 ;
        RECT 79.215 150.825 79.385 150.995 ;
        RECT 79.675 150.825 79.845 150.995 ;
        RECT 80.135 150.825 80.305 150.995 ;
        RECT 80.595 150.825 80.765 150.995 ;
        RECT 81.055 150.825 81.225 150.995 ;
        RECT 81.515 150.825 81.685 150.995 ;
        RECT 81.975 150.825 82.145 150.995 ;
        RECT 82.435 150.825 82.605 150.995 ;
        RECT 82.895 150.825 83.065 150.995 ;
        RECT 83.355 150.825 83.525 150.995 ;
        RECT 83.815 150.825 83.985 150.995 ;
        RECT 84.275 150.825 84.445 150.995 ;
        RECT 84.735 150.825 84.905 150.995 ;
        RECT 85.195 150.825 85.365 150.995 ;
        RECT 85.655 150.825 85.825 150.995 ;
        RECT 86.115 150.825 86.285 150.995 ;
        RECT 86.575 150.825 86.745 150.995 ;
        RECT 87.035 150.825 87.205 150.995 ;
        RECT 87.495 150.825 87.665 150.995 ;
        RECT 87.955 150.825 88.125 150.995 ;
        RECT 88.415 150.825 88.585 150.995 ;
        RECT 88.875 150.825 89.045 150.995 ;
        RECT 89.335 150.825 89.505 150.995 ;
        RECT 89.795 150.825 89.965 150.995 ;
        RECT 90.255 150.825 90.425 150.995 ;
        RECT 90.715 150.825 90.885 150.995 ;
        RECT 91.175 150.825 91.345 150.995 ;
        RECT 91.635 150.825 91.805 150.995 ;
        RECT 92.095 150.825 92.265 150.995 ;
        RECT 92.555 150.825 92.725 150.995 ;
        RECT 93.015 150.825 93.185 150.995 ;
        RECT 93.475 150.825 93.645 150.995 ;
        RECT 93.935 150.825 94.105 150.995 ;
        RECT 94.395 150.825 94.565 150.995 ;
        RECT 94.855 150.825 95.025 150.995 ;
        RECT 95.315 150.825 95.485 150.995 ;
        RECT 95.775 150.825 95.945 150.995 ;
        RECT 96.235 150.825 96.405 150.995 ;
        RECT 96.695 150.825 96.865 150.995 ;
        RECT 97.155 150.825 97.325 150.995 ;
        RECT 97.615 150.825 97.785 150.995 ;
        RECT 98.075 150.825 98.245 150.995 ;
        RECT 98.535 150.825 98.705 150.995 ;
        RECT 98.995 150.825 99.165 150.995 ;
        RECT 99.455 150.825 99.625 150.995 ;
        RECT 99.915 150.825 100.085 150.995 ;
        RECT 100.375 150.825 100.545 150.995 ;
        RECT 100.835 150.825 101.005 150.995 ;
        RECT 101.295 150.825 101.465 150.995 ;
        RECT 101.755 150.825 101.925 150.995 ;
        RECT 102.215 150.825 102.385 150.995 ;
        RECT 102.675 150.825 102.845 150.995 ;
        RECT 103.135 150.825 103.305 150.995 ;
        RECT 103.595 150.825 103.765 150.995 ;
        RECT 104.055 150.825 104.225 150.995 ;
        RECT 104.515 150.825 104.685 150.995 ;
        RECT 104.975 150.825 105.145 150.995 ;
        RECT 105.435 150.825 105.605 150.995 ;
        RECT 105.895 150.825 106.065 150.995 ;
        RECT 106.355 150.825 106.525 150.995 ;
        RECT 106.815 150.825 106.985 150.995 ;
        RECT 107.275 150.825 107.445 150.995 ;
        RECT 107.735 150.825 107.905 150.995 ;
        RECT 108.195 150.825 108.365 150.995 ;
        RECT 108.655 150.825 108.825 150.995 ;
        RECT 109.115 150.825 109.285 150.995 ;
        RECT 109.575 150.825 109.745 150.995 ;
        RECT 110.035 150.825 110.205 150.995 ;
        RECT 110.495 150.825 110.665 150.995 ;
        RECT 110.955 150.825 111.125 150.995 ;
        RECT 111.415 150.825 111.585 150.995 ;
        RECT 111.875 150.825 112.045 150.995 ;
        RECT 112.335 150.825 112.505 150.995 ;
        RECT 112.795 150.825 112.965 150.995 ;
        RECT 113.255 150.825 113.425 150.995 ;
        RECT 113.715 150.825 113.885 150.995 ;
        RECT 114.175 150.825 114.345 150.995 ;
        RECT 114.635 150.825 114.805 150.995 ;
        RECT 115.095 150.825 115.265 150.995 ;
        RECT 115.555 150.825 115.725 150.995 ;
        RECT 116.015 150.825 116.185 150.995 ;
        RECT 116.475 150.825 116.645 150.995 ;
        RECT 116.935 150.825 117.105 150.995 ;
        RECT 117.395 150.825 117.565 150.995 ;
        RECT 117.855 150.825 118.025 150.995 ;
        RECT 118.315 150.825 118.485 150.995 ;
        RECT 118.775 150.825 118.945 150.995 ;
        RECT 119.235 150.825 119.405 150.995 ;
        RECT 21.130 150.320 21.300 150.490 ;
        RECT 81.055 150.315 81.225 150.485 ;
        RECT 81.975 149.295 82.145 149.465 ;
        RECT 84.735 149.635 84.905 149.805 ;
        RECT 85.200 149.295 85.370 149.465 ;
        RECT 85.605 149.975 85.775 150.145 ;
        RECT 86.115 148.955 86.285 149.125 ;
        RECT 87.495 149.975 87.665 150.145 ;
        RECT 87.035 149.295 87.205 149.465 ;
        RECT 90.615 149.975 90.785 150.145 ;
        RECT 88.755 148.955 88.925 149.125 ;
        RECT 90.615 149.295 90.785 149.465 ;
        RECT 93.475 150.315 93.645 150.485 ;
        RECT 91.695 149.270 91.865 149.440 ;
        RECT 91.995 148.955 92.165 149.125 ;
        RECT 104.515 149.295 104.685 149.465 ;
        RECT 105.435 148.615 105.605 148.785 ;
        RECT 105.895 150.315 106.065 150.485 ;
        RECT 106.815 149.295 106.985 149.465 ;
        RECT 107.275 149.295 107.445 149.465 ;
        RECT 107.735 149.975 107.905 150.145 ;
        RECT 108.195 149.295 108.365 149.465 ;
        RECT 110.495 149.295 110.665 149.465 ;
        RECT 114.635 150.315 114.805 150.485 ;
        RECT 113.255 149.635 113.425 149.805 ;
        RECT 117.855 149.635 118.025 149.805 ;
        RECT 71.395 148.105 71.565 148.275 ;
        RECT 71.855 148.105 72.025 148.275 ;
        RECT 72.315 148.105 72.485 148.275 ;
        RECT 72.775 148.105 72.945 148.275 ;
        RECT 73.235 148.105 73.405 148.275 ;
        RECT 73.695 148.105 73.865 148.275 ;
        RECT 74.155 148.105 74.325 148.275 ;
        RECT 74.615 148.105 74.785 148.275 ;
        RECT 75.075 148.105 75.245 148.275 ;
        RECT 75.535 148.105 75.705 148.275 ;
        RECT 75.995 148.105 76.165 148.275 ;
        RECT 76.455 148.105 76.625 148.275 ;
        RECT 76.915 148.105 77.085 148.275 ;
        RECT 77.375 148.105 77.545 148.275 ;
        RECT 77.835 148.105 78.005 148.275 ;
        RECT 78.295 148.105 78.465 148.275 ;
        RECT 78.755 148.105 78.925 148.275 ;
        RECT 79.215 148.105 79.385 148.275 ;
        RECT 79.675 148.105 79.845 148.275 ;
        RECT 80.135 148.105 80.305 148.275 ;
        RECT 80.595 148.105 80.765 148.275 ;
        RECT 81.055 148.105 81.225 148.275 ;
        RECT 81.515 148.105 81.685 148.275 ;
        RECT 81.975 148.105 82.145 148.275 ;
        RECT 82.435 148.105 82.605 148.275 ;
        RECT 82.895 148.105 83.065 148.275 ;
        RECT 83.355 148.105 83.525 148.275 ;
        RECT 83.815 148.105 83.985 148.275 ;
        RECT 84.275 148.105 84.445 148.275 ;
        RECT 84.735 148.105 84.905 148.275 ;
        RECT 85.195 148.105 85.365 148.275 ;
        RECT 85.655 148.105 85.825 148.275 ;
        RECT 86.115 148.105 86.285 148.275 ;
        RECT 86.575 148.105 86.745 148.275 ;
        RECT 87.035 148.105 87.205 148.275 ;
        RECT 87.495 148.105 87.665 148.275 ;
        RECT 87.955 148.105 88.125 148.275 ;
        RECT 88.415 148.105 88.585 148.275 ;
        RECT 88.875 148.105 89.045 148.275 ;
        RECT 89.335 148.105 89.505 148.275 ;
        RECT 89.795 148.105 89.965 148.275 ;
        RECT 90.255 148.105 90.425 148.275 ;
        RECT 90.715 148.105 90.885 148.275 ;
        RECT 91.175 148.105 91.345 148.275 ;
        RECT 91.635 148.105 91.805 148.275 ;
        RECT 92.095 148.105 92.265 148.275 ;
        RECT 92.555 148.105 92.725 148.275 ;
        RECT 93.015 148.105 93.185 148.275 ;
        RECT 93.475 148.105 93.645 148.275 ;
        RECT 93.935 148.105 94.105 148.275 ;
        RECT 94.395 148.105 94.565 148.275 ;
        RECT 94.855 148.105 95.025 148.275 ;
        RECT 95.315 148.105 95.485 148.275 ;
        RECT 95.775 148.105 95.945 148.275 ;
        RECT 96.235 148.105 96.405 148.275 ;
        RECT 96.695 148.105 96.865 148.275 ;
        RECT 97.155 148.105 97.325 148.275 ;
        RECT 97.615 148.105 97.785 148.275 ;
        RECT 98.075 148.105 98.245 148.275 ;
        RECT 98.535 148.105 98.705 148.275 ;
        RECT 98.995 148.105 99.165 148.275 ;
        RECT 99.455 148.105 99.625 148.275 ;
        RECT 99.915 148.105 100.085 148.275 ;
        RECT 100.375 148.105 100.545 148.275 ;
        RECT 100.835 148.105 101.005 148.275 ;
        RECT 101.295 148.105 101.465 148.275 ;
        RECT 101.755 148.105 101.925 148.275 ;
        RECT 102.215 148.105 102.385 148.275 ;
        RECT 102.675 148.105 102.845 148.275 ;
        RECT 103.135 148.105 103.305 148.275 ;
        RECT 103.595 148.105 103.765 148.275 ;
        RECT 104.055 148.105 104.225 148.275 ;
        RECT 104.515 148.105 104.685 148.275 ;
        RECT 104.975 148.105 105.145 148.275 ;
        RECT 105.435 148.105 105.605 148.275 ;
        RECT 105.895 148.105 106.065 148.275 ;
        RECT 106.355 148.105 106.525 148.275 ;
        RECT 106.815 148.105 106.985 148.275 ;
        RECT 107.275 148.105 107.445 148.275 ;
        RECT 107.735 148.105 107.905 148.275 ;
        RECT 108.195 148.105 108.365 148.275 ;
        RECT 108.655 148.105 108.825 148.275 ;
        RECT 109.115 148.105 109.285 148.275 ;
        RECT 109.575 148.105 109.745 148.275 ;
        RECT 110.035 148.105 110.205 148.275 ;
        RECT 110.495 148.105 110.665 148.275 ;
        RECT 110.955 148.105 111.125 148.275 ;
        RECT 111.415 148.105 111.585 148.275 ;
        RECT 111.875 148.105 112.045 148.275 ;
        RECT 112.335 148.105 112.505 148.275 ;
        RECT 112.795 148.105 112.965 148.275 ;
        RECT 113.255 148.105 113.425 148.275 ;
        RECT 113.715 148.105 113.885 148.275 ;
        RECT 114.175 148.105 114.345 148.275 ;
        RECT 114.635 148.105 114.805 148.275 ;
        RECT 115.095 148.105 115.265 148.275 ;
        RECT 115.555 148.105 115.725 148.275 ;
        RECT 116.015 148.105 116.185 148.275 ;
        RECT 116.475 148.105 116.645 148.275 ;
        RECT 116.935 148.105 117.105 148.275 ;
        RECT 117.395 148.105 117.565 148.275 ;
        RECT 117.855 148.105 118.025 148.275 ;
        RECT 118.315 148.105 118.485 148.275 ;
        RECT 118.775 148.105 118.945 148.275 ;
        RECT 119.235 148.105 119.405 148.275 ;
        RECT 12.655 135.580 12.825 136.460 ;
        RECT 13.095 135.580 13.265 136.460 ;
        RECT 12.650 132.605 12.840 134.590 ;
        RECT 17.210 136.440 17.380 136.610 ;
        RECT 18.000 135.475 18.170 135.645 ;
        RECT 17.780 134.345 17.950 135.225 ;
        RECT 18.220 134.345 18.390 135.225 ;
        RECT 20.030 135.475 20.200 135.645 ;
        RECT 18.000 133.925 18.170 134.095 ;
        RECT 19.810 134.345 19.980 135.225 ;
        RECT 20.250 134.345 20.420 135.225 ;
        RECT 20.030 133.925 20.200 134.095 ;
        RECT 22.060 135.475 22.230 135.645 ;
        RECT 21.840 134.345 22.010 135.225 ;
        RECT 22.280 134.345 22.450 135.225 ;
        RECT 22.060 133.925 22.230 134.095 ;
        RECT 24.090 135.485 24.260 135.655 ;
        RECT 23.870 134.355 24.040 135.235 ;
        RECT 24.310 134.355 24.480 135.235 ;
        RECT 24.090 133.935 24.260 134.105 ;
        RECT 26.110 135.485 26.280 135.655 ;
        RECT 25.890 134.355 26.060 135.235 ;
        RECT 26.330 134.355 26.500 135.235 ;
        RECT 28.135 135.480 28.305 135.650 ;
        RECT 26.110 133.935 26.280 134.105 ;
        RECT 27.915 134.350 28.085 135.230 ;
        RECT 28.355 134.350 28.525 135.230 ;
        RECT 28.135 133.930 28.305 134.100 ;
        RECT 12.650 129.950 12.840 131.935 ;
        RECT 17.495 115.035 17.670 115.220 ;
        RECT 20.500 115.055 20.670 115.230 ;
        RECT 14.650 109.065 15.280 109.635 ;
        RECT 18.740 113.255 18.910 114.135 ;
        RECT 19.180 113.255 19.350 114.135 ;
        RECT 19.620 113.255 19.790 114.135 ;
        RECT 20.250 113.255 20.420 114.135 ;
        RECT 20.690 113.255 20.860 114.135 ;
        RECT 21.130 113.255 21.300 114.135 ;
        RECT 20.910 112.350 21.080 112.520 ;
        RECT 12.435 97.610 12.605 98.490 ;
        RECT 12.875 97.610 13.045 98.490 ;
        RECT 12.430 94.635 12.620 96.620 ;
        RECT 16.990 98.470 17.160 98.640 ;
        RECT 17.780 97.505 17.950 97.675 ;
        RECT 17.560 96.375 17.730 97.255 ;
        RECT 18.000 96.375 18.170 97.255 ;
        RECT 19.810 97.505 19.980 97.675 ;
        RECT 17.780 95.955 17.950 96.125 ;
        RECT 19.590 96.375 19.760 97.255 ;
        RECT 20.030 96.375 20.200 97.255 ;
        RECT 19.810 95.955 19.980 96.125 ;
        RECT 21.840 97.505 22.010 97.675 ;
        RECT 21.620 96.375 21.790 97.255 ;
        RECT 22.060 96.375 22.230 97.255 ;
        RECT 21.840 95.955 22.010 96.125 ;
        RECT 23.870 97.515 24.040 97.685 ;
        RECT 23.650 96.385 23.820 97.265 ;
        RECT 24.090 96.385 24.260 97.265 ;
        RECT 23.870 95.965 24.040 96.135 ;
        RECT 25.890 97.515 26.060 97.685 ;
        RECT 25.670 96.385 25.840 97.265 ;
        RECT 26.110 96.385 26.280 97.265 ;
        RECT 27.915 97.510 28.085 97.680 ;
        RECT 25.890 95.965 26.060 96.135 ;
        RECT 27.695 96.380 27.865 97.260 ;
        RECT 28.135 96.380 28.305 97.260 ;
        RECT 27.915 95.960 28.085 96.130 ;
        RECT 12.430 91.980 12.620 93.965 ;
        RECT 91.205 88.855 91.375 89.025 ;
        RECT 91.665 88.855 91.835 89.025 ;
        RECT 92.125 88.855 92.295 89.025 ;
        RECT 92.585 88.855 92.755 89.025 ;
        RECT 93.045 88.855 93.215 89.025 ;
        RECT 93.505 88.855 93.675 89.025 ;
        RECT 93.965 88.855 94.135 89.025 ;
        RECT 94.425 88.855 94.595 89.025 ;
        RECT 94.885 88.855 95.055 89.025 ;
        RECT 95.345 88.855 95.515 89.025 ;
        RECT 95.805 88.855 95.975 89.025 ;
        RECT 96.265 88.855 96.435 89.025 ;
        RECT 96.725 88.855 96.895 89.025 ;
        RECT 97.185 88.855 97.355 89.025 ;
        RECT 97.645 88.855 97.815 89.025 ;
        RECT 98.105 88.855 98.275 89.025 ;
        RECT 98.565 88.855 98.735 89.025 ;
        RECT 99.025 88.855 99.195 89.025 ;
        RECT 99.485 88.855 99.655 89.025 ;
        RECT 99.945 88.855 100.115 89.025 ;
        RECT 100.405 88.855 100.575 89.025 ;
        RECT 100.865 88.855 101.035 89.025 ;
        RECT 101.325 88.855 101.495 89.025 ;
        RECT 101.785 88.855 101.955 89.025 ;
        RECT 102.245 88.855 102.415 89.025 ;
        RECT 102.705 88.855 102.875 89.025 ;
        RECT 103.165 88.855 103.335 89.025 ;
        RECT 103.625 88.855 103.795 89.025 ;
        RECT 104.085 88.855 104.255 89.025 ;
        RECT 104.545 88.855 104.715 89.025 ;
        RECT 105.005 88.855 105.175 89.025 ;
        RECT 105.465 88.855 105.635 89.025 ;
        RECT 105.925 88.855 106.095 89.025 ;
        RECT 106.385 88.855 106.555 89.025 ;
        RECT 106.845 88.855 107.015 89.025 ;
        RECT 107.305 88.855 107.475 89.025 ;
        RECT 107.765 88.855 107.935 89.025 ;
        RECT 108.225 88.855 108.395 89.025 ;
        RECT 108.685 88.855 108.855 89.025 ;
        RECT 109.145 88.855 109.315 89.025 ;
        RECT 109.605 88.855 109.775 89.025 ;
        RECT 110.065 88.855 110.235 89.025 ;
        RECT 110.525 88.855 110.695 89.025 ;
        RECT 110.985 88.855 111.155 89.025 ;
        RECT 111.445 88.855 111.615 89.025 ;
        RECT 111.905 88.855 112.075 89.025 ;
        RECT 112.365 88.855 112.535 89.025 ;
        RECT 112.825 88.855 112.995 89.025 ;
        RECT 113.285 88.855 113.455 89.025 ;
        RECT 113.745 88.855 113.915 89.025 ;
        RECT 114.205 88.855 114.375 89.025 ;
        RECT 114.665 88.855 114.835 89.025 ;
        RECT 115.125 88.855 115.295 89.025 ;
        RECT 115.585 88.855 115.755 89.025 ;
        RECT 116.045 88.855 116.215 89.025 ;
        RECT 116.505 88.855 116.675 89.025 ;
        RECT 116.965 88.855 117.135 89.025 ;
        RECT 117.425 88.855 117.595 89.025 ;
        RECT 117.885 88.855 118.055 89.025 ;
        RECT 118.345 88.855 118.515 89.025 ;
        RECT 118.805 88.855 118.975 89.025 ;
        RECT 119.265 88.855 119.435 89.025 ;
        RECT 119.725 88.855 119.895 89.025 ;
        RECT 120.185 88.855 120.355 89.025 ;
        RECT 120.645 88.855 120.815 89.025 ;
        RECT 121.105 88.855 121.275 89.025 ;
        RECT 121.565 88.855 121.735 89.025 ;
        RECT 122.025 88.855 122.195 89.025 ;
        RECT 122.485 88.855 122.655 89.025 ;
        RECT 122.945 88.855 123.115 89.025 ;
        RECT 123.405 88.855 123.575 89.025 ;
        RECT 123.865 88.855 124.035 89.025 ;
        RECT 124.325 88.855 124.495 89.025 ;
        RECT 124.785 88.855 124.955 89.025 ;
        RECT 125.245 88.855 125.415 89.025 ;
        RECT 125.705 88.855 125.875 89.025 ;
        RECT 126.165 88.855 126.335 89.025 ;
        RECT 126.625 88.855 126.795 89.025 ;
        RECT 127.085 88.855 127.255 89.025 ;
        RECT 127.545 88.855 127.715 89.025 ;
        RECT 128.005 88.855 128.175 89.025 ;
        RECT 128.465 88.855 128.635 89.025 ;
        RECT 128.925 88.855 129.095 89.025 ;
        RECT 129.385 88.855 129.555 89.025 ;
        RECT 129.845 88.855 130.015 89.025 ;
        RECT 130.305 88.855 130.475 89.025 ;
        RECT 130.765 88.855 130.935 89.025 ;
        RECT 131.225 88.855 131.395 89.025 ;
        RECT 131.685 88.855 131.855 89.025 ;
        RECT 132.145 88.855 132.315 89.025 ;
        RECT 132.605 88.855 132.775 89.025 ;
        RECT 133.065 88.855 133.235 89.025 ;
        RECT 133.525 88.855 133.695 89.025 ;
        RECT 133.985 88.855 134.155 89.025 ;
        RECT 134.445 88.855 134.615 89.025 ;
        RECT 134.905 88.855 135.075 89.025 ;
        RECT 135.365 88.855 135.535 89.025 ;
        RECT 135.825 88.855 135.995 89.025 ;
        RECT 136.285 88.855 136.455 89.025 ;
        RECT 136.745 88.855 136.915 89.025 ;
        RECT 137.205 88.855 137.375 89.025 ;
        RECT 137.665 88.855 137.835 89.025 ;
        RECT 138.125 88.855 138.295 89.025 ;
        RECT 138.585 88.855 138.755 89.025 ;
        RECT 139.045 88.855 139.215 89.025 ;
        RECT 139.505 88.855 139.675 89.025 ;
        RECT 139.965 88.855 140.135 89.025 ;
        RECT 140.425 88.855 140.595 89.025 ;
        RECT 140.885 88.855 141.055 89.025 ;
        RECT 141.345 88.855 141.515 89.025 ;
        RECT 141.805 88.855 141.975 89.025 ;
        RECT 142.265 88.855 142.435 89.025 ;
        RECT 142.725 88.855 142.895 89.025 ;
        RECT 143.185 88.855 143.355 89.025 ;
        RECT 143.645 88.855 143.815 89.025 ;
        RECT 144.105 88.855 144.275 89.025 ;
        RECT 144.565 88.855 144.735 89.025 ;
        RECT 145.025 88.855 145.195 89.025 ;
        RECT 145.485 88.855 145.655 89.025 ;
        RECT 145.945 88.855 146.115 89.025 ;
        RECT 146.405 88.855 146.575 89.025 ;
        RECT 146.865 88.855 147.035 89.025 ;
        RECT 147.325 88.855 147.495 89.025 ;
        RECT 147.785 88.855 147.955 89.025 ;
        RECT 148.245 88.855 148.415 89.025 ;
        RECT 148.705 88.855 148.875 89.025 ;
        RECT 149.165 88.855 149.335 89.025 ;
        RECT 149.625 88.855 149.795 89.025 ;
        RECT 150.085 88.855 150.255 89.025 ;
        RECT 150.545 88.855 150.715 89.025 ;
        RECT 151.005 88.855 151.175 89.025 ;
        RECT 151.465 88.855 151.635 89.025 ;
        RECT 151.925 88.855 152.095 89.025 ;
        RECT 105.005 88.345 105.175 88.515 ;
        RECT 106.385 87.665 106.555 87.835 ;
        RECT 140.885 88.345 141.055 88.515 ;
        RECT 140.425 87.665 140.595 87.835 ;
        RECT 150.085 88.005 150.255 88.175 ;
        RECT 149.165 86.985 149.335 87.155 ;
        RECT 91.205 86.135 91.375 86.305 ;
        RECT 91.665 86.135 91.835 86.305 ;
        RECT 92.125 86.135 92.295 86.305 ;
        RECT 92.585 86.135 92.755 86.305 ;
        RECT 93.045 86.135 93.215 86.305 ;
        RECT 93.505 86.135 93.675 86.305 ;
        RECT 93.965 86.135 94.135 86.305 ;
        RECT 94.425 86.135 94.595 86.305 ;
        RECT 94.885 86.135 95.055 86.305 ;
        RECT 95.345 86.135 95.515 86.305 ;
        RECT 95.805 86.135 95.975 86.305 ;
        RECT 96.265 86.135 96.435 86.305 ;
        RECT 96.725 86.135 96.895 86.305 ;
        RECT 97.185 86.135 97.355 86.305 ;
        RECT 97.645 86.135 97.815 86.305 ;
        RECT 98.105 86.135 98.275 86.305 ;
        RECT 98.565 86.135 98.735 86.305 ;
        RECT 99.025 86.135 99.195 86.305 ;
        RECT 99.485 86.135 99.655 86.305 ;
        RECT 99.945 86.135 100.115 86.305 ;
        RECT 100.405 86.135 100.575 86.305 ;
        RECT 100.865 86.135 101.035 86.305 ;
        RECT 101.325 86.135 101.495 86.305 ;
        RECT 101.785 86.135 101.955 86.305 ;
        RECT 102.245 86.135 102.415 86.305 ;
        RECT 102.705 86.135 102.875 86.305 ;
        RECT 103.165 86.135 103.335 86.305 ;
        RECT 103.625 86.135 103.795 86.305 ;
        RECT 104.085 86.135 104.255 86.305 ;
        RECT 104.545 86.135 104.715 86.305 ;
        RECT 105.005 86.135 105.175 86.305 ;
        RECT 105.465 86.135 105.635 86.305 ;
        RECT 105.925 86.135 106.095 86.305 ;
        RECT 106.385 86.135 106.555 86.305 ;
        RECT 106.845 86.135 107.015 86.305 ;
        RECT 107.305 86.135 107.475 86.305 ;
        RECT 107.765 86.135 107.935 86.305 ;
        RECT 108.225 86.135 108.395 86.305 ;
        RECT 108.685 86.135 108.855 86.305 ;
        RECT 109.145 86.135 109.315 86.305 ;
        RECT 109.605 86.135 109.775 86.305 ;
        RECT 110.065 86.135 110.235 86.305 ;
        RECT 110.525 86.135 110.695 86.305 ;
        RECT 110.985 86.135 111.155 86.305 ;
        RECT 111.445 86.135 111.615 86.305 ;
        RECT 111.905 86.135 112.075 86.305 ;
        RECT 112.365 86.135 112.535 86.305 ;
        RECT 112.825 86.135 112.995 86.305 ;
        RECT 113.285 86.135 113.455 86.305 ;
        RECT 113.745 86.135 113.915 86.305 ;
        RECT 114.205 86.135 114.375 86.305 ;
        RECT 114.665 86.135 114.835 86.305 ;
        RECT 115.125 86.135 115.295 86.305 ;
        RECT 115.585 86.135 115.755 86.305 ;
        RECT 116.045 86.135 116.215 86.305 ;
        RECT 116.505 86.135 116.675 86.305 ;
        RECT 116.965 86.135 117.135 86.305 ;
        RECT 117.425 86.135 117.595 86.305 ;
        RECT 117.885 86.135 118.055 86.305 ;
        RECT 118.345 86.135 118.515 86.305 ;
        RECT 118.805 86.135 118.975 86.305 ;
        RECT 119.265 86.135 119.435 86.305 ;
        RECT 119.725 86.135 119.895 86.305 ;
        RECT 120.185 86.135 120.355 86.305 ;
        RECT 120.645 86.135 120.815 86.305 ;
        RECT 121.105 86.135 121.275 86.305 ;
        RECT 121.565 86.135 121.735 86.305 ;
        RECT 122.025 86.135 122.195 86.305 ;
        RECT 122.485 86.135 122.655 86.305 ;
        RECT 122.945 86.135 123.115 86.305 ;
        RECT 123.405 86.135 123.575 86.305 ;
        RECT 123.865 86.135 124.035 86.305 ;
        RECT 124.325 86.135 124.495 86.305 ;
        RECT 124.785 86.135 124.955 86.305 ;
        RECT 125.245 86.135 125.415 86.305 ;
        RECT 125.705 86.135 125.875 86.305 ;
        RECT 126.165 86.135 126.335 86.305 ;
        RECT 126.625 86.135 126.795 86.305 ;
        RECT 127.085 86.135 127.255 86.305 ;
        RECT 127.545 86.135 127.715 86.305 ;
        RECT 128.005 86.135 128.175 86.305 ;
        RECT 128.465 86.135 128.635 86.305 ;
        RECT 128.925 86.135 129.095 86.305 ;
        RECT 129.385 86.135 129.555 86.305 ;
        RECT 129.845 86.135 130.015 86.305 ;
        RECT 130.305 86.135 130.475 86.305 ;
        RECT 130.765 86.135 130.935 86.305 ;
        RECT 131.225 86.135 131.395 86.305 ;
        RECT 131.685 86.135 131.855 86.305 ;
        RECT 132.145 86.135 132.315 86.305 ;
        RECT 132.605 86.135 132.775 86.305 ;
        RECT 133.065 86.135 133.235 86.305 ;
        RECT 133.525 86.135 133.695 86.305 ;
        RECT 133.985 86.135 134.155 86.305 ;
        RECT 134.445 86.135 134.615 86.305 ;
        RECT 134.905 86.135 135.075 86.305 ;
        RECT 135.365 86.135 135.535 86.305 ;
        RECT 135.825 86.135 135.995 86.305 ;
        RECT 136.285 86.135 136.455 86.305 ;
        RECT 136.745 86.135 136.915 86.305 ;
        RECT 137.205 86.135 137.375 86.305 ;
        RECT 137.665 86.135 137.835 86.305 ;
        RECT 138.125 86.135 138.295 86.305 ;
        RECT 138.585 86.135 138.755 86.305 ;
        RECT 139.045 86.135 139.215 86.305 ;
        RECT 139.505 86.135 139.675 86.305 ;
        RECT 139.965 86.135 140.135 86.305 ;
        RECT 140.425 86.135 140.595 86.305 ;
        RECT 140.885 86.135 141.055 86.305 ;
        RECT 141.345 86.135 141.515 86.305 ;
        RECT 141.805 86.135 141.975 86.305 ;
        RECT 142.265 86.135 142.435 86.305 ;
        RECT 142.725 86.135 142.895 86.305 ;
        RECT 143.185 86.135 143.355 86.305 ;
        RECT 143.645 86.135 143.815 86.305 ;
        RECT 144.105 86.135 144.275 86.305 ;
        RECT 144.565 86.135 144.735 86.305 ;
        RECT 145.025 86.135 145.195 86.305 ;
        RECT 145.485 86.135 145.655 86.305 ;
        RECT 145.945 86.135 146.115 86.305 ;
        RECT 146.405 86.135 146.575 86.305 ;
        RECT 146.865 86.135 147.035 86.305 ;
        RECT 147.325 86.135 147.495 86.305 ;
        RECT 147.785 86.135 147.955 86.305 ;
        RECT 148.245 86.135 148.415 86.305 ;
        RECT 148.705 86.135 148.875 86.305 ;
        RECT 149.165 86.135 149.335 86.305 ;
        RECT 149.625 86.135 149.795 86.305 ;
        RECT 150.085 86.135 150.255 86.305 ;
        RECT 150.545 86.135 150.715 86.305 ;
        RECT 151.005 86.135 151.175 86.305 ;
        RECT 151.465 86.135 151.635 86.305 ;
        RECT 151.925 86.135 152.095 86.305 ;
        RECT 122.025 84.605 122.195 84.775 ;
        RECT 122.945 84.605 123.115 84.775 ;
        RECT 122.945 83.925 123.115 84.095 ;
        RECT 126.165 84.605 126.335 84.775 ;
        RECT 130.305 84.605 130.475 84.775 ;
        RECT 131.225 84.605 131.395 84.775 ;
        RECT 132.145 84.605 132.315 84.775 ;
        RECT 125.245 83.925 125.415 84.095 ;
        RECT 133.985 84.605 134.155 84.775 ;
        RECT 134.905 83.925 135.075 84.095 ;
        RECT 136.745 84.945 136.915 85.115 ;
        RECT 137.210 84.605 137.380 84.775 ;
        RECT 137.615 85.285 137.785 85.455 ;
        RECT 138.125 84.265 138.295 84.435 ;
        RECT 139.505 85.285 139.675 85.455 ;
        RECT 139.045 84.605 139.215 84.775 ;
        RECT 142.625 85.285 142.795 85.455 ;
        RECT 140.765 84.265 140.935 84.435 ;
        RECT 142.625 84.605 142.795 84.775 ;
        RECT 143.705 84.580 143.875 84.750 ;
        RECT 144.005 84.265 144.175 84.435 ;
        RECT 145.485 83.925 145.655 84.095 ;
        RECT 91.205 83.415 91.375 83.585 ;
        RECT 91.665 83.415 91.835 83.585 ;
        RECT 92.125 83.415 92.295 83.585 ;
        RECT 92.585 83.415 92.755 83.585 ;
        RECT 93.045 83.415 93.215 83.585 ;
        RECT 93.505 83.415 93.675 83.585 ;
        RECT 93.965 83.415 94.135 83.585 ;
        RECT 94.425 83.415 94.595 83.585 ;
        RECT 94.885 83.415 95.055 83.585 ;
        RECT 95.345 83.415 95.515 83.585 ;
        RECT 95.805 83.415 95.975 83.585 ;
        RECT 96.265 83.415 96.435 83.585 ;
        RECT 96.725 83.415 96.895 83.585 ;
        RECT 97.185 83.415 97.355 83.585 ;
        RECT 97.645 83.415 97.815 83.585 ;
        RECT 98.105 83.415 98.275 83.585 ;
        RECT 98.565 83.415 98.735 83.585 ;
        RECT 99.025 83.415 99.195 83.585 ;
        RECT 99.485 83.415 99.655 83.585 ;
        RECT 99.945 83.415 100.115 83.585 ;
        RECT 100.405 83.415 100.575 83.585 ;
        RECT 100.865 83.415 101.035 83.585 ;
        RECT 101.325 83.415 101.495 83.585 ;
        RECT 101.785 83.415 101.955 83.585 ;
        RECT 102.245 83.415 102.415 83.585 ;
        RECT 102.705 83.415 102.875 83.585 ;
        RECT 103.165 83.415 103.335 83.585 ;
        RECT 103.625 83.415 103.795 83.585 ;
        RECT 104.085 83.415 104.255 83.585 ;
        RECT 104.545 83.415 104.715 83.585 ;
        RECT 105.005 83.415 105.175 83.585 ;
        RECT 105.465 83.415 105.635 83.585 ;
        RECT 105.925 83.415 106.095 83.585 ;
        RECT 106.385 83.415 106.555 83.585 ;
        RECT 106.845 83.415 107.015 83.585 ;
        RECT 107.305 83.415 107.475 83.585 ;
        RECT 107.765 83.415 107.935 83.585 ;
        RECT 108.225 83.415 108.395 83.585 ;
        RECT 108.685 83.415 108.855 83.585 ;
        RECT 109.145 83.415 109.315 83.585 ;
        RECT 109.605 83.415 109.775 83.585 ;
        RECT 110.065 83.415 110.235 83.585 ;
        RECT 110.525 83.415 110.695 83.585 ;
        RECT 110.985 83.415 111.155 83.585 ;
        RECT 111.445 83.415 111.615 83.585 ;
        RECT 111.905 83.415 112.075 83.585 ;
        RECT 112.365 83.415 112.535 83.585 ;
        RECT 112.825 83.415 112.995 83.585 ;
        RECT 113.285 83.415 113.455 83.585 ;
        RECT 113.745 83.415 113.915 83.585 ;
        RECT 114.205 83.415 114.375 83.585 ;
        RECT 114.665 83.415 114.835 83.585 ;
        RECT 115.125 83.415 115.295 83.585 ;
        RECT 115.585 83.415 115.755 83.585 ;
        RECT 116.045 83.415 116.215 83.585 ;
        RECT 116.505 83.415 116.675 83.585 ;
        RECT 116.965 83.415 117.135 83.585 ;
        RECT 117.425 83.415 117.595 83.585 ;
        RECT 117.885 83.415 118.055 83.585 ;
        RECT 118.345 83.415 118.515 83.585 ;
        RECT 118.805 83.415 118.975 83.585 ;
        RECT 119.265 83.415 119.435 83.585 ;
        RECT 119.725 83.415 119.895 83.585 ;
        RECT 120.185 83.415 120.355 83.585 ;
        RECT 120.645 83.415 120.815 83.585 ;
        RECT 121.105 83.415 121.275 83.585 ;
        RECT 121.565 83.415 121.735 83.585 ;
        RECT 122.025 83.415 122.195 83.585 ;
        RECT 122.485 83.415 122.655 83.585 ;
        RECT 122.945 83.415 123.115 83.585 ;
        RECT 123.405 83.415 123.575 83.585 ;
        RECT 123.865 83.415 124.035 83.585 ;
        RECT 124.325 83.415 124.495 83.585 ;
        RECT 124.785 83.415 124.955 83.585 ;
        RECT 125.245 83.415 125.415 83.585 ;
        RECT 125.705 83.415 125.875 83.585 ;
        RECT 126.165 83.415 126.335 83.585 ;
        RECT 126.625 83.415 126.795 83.585 ;
        RECT 127.085 83.415 127.255 83.585 ;
        RECT 127.545 83.415 127.715 83.585 ;
        RECT 128.005 83.415 128.175 83.585 ;
        RECT 128.465 83.415 128.635 83.585 ;
        RECT 128.925 83.415 129.095 83.585 ;
        RECT 129.385 83.415 129.555 83.585 ;
        RECT 129.845 83.415 130.015 83.585 ;
        RECT 130.305 83.415 130.475 83.585 ;
        RECT 130.765 83.415 130.935 83.585 ;
        RECT 131.225 83.415 131.395 83.585 ;
        RECT 131.685 83.415 131.855 83.585 ;
        RECT 132.145 83.415 132.315 83.585 ;
        RECT 132.605 83.415 132.775 83.585 ;
        RECT 133.065 83.415 133.235 83.585 ;
        RECT 133.525 83.415 133.695 83.585 ;
        RECT 133.985 83.415 134.155 83.585 ;
        RECT 134.445 83.415 134.615 83.585 ;
        RECT 134.905 83.415 135.075 83.585 ;
        RECT 135.365 83.415 135.535 83.585 ;
        RECT 135.825 83.415 135.995 83.585 ;
        RECT 136.285 83.415 136.455 83.585 ;
        RECT 136.745 83.415 136.915 83.585 ;
        RECT 137.205 83.415 137.375 83.585 ;
        RECT 137.665 83.415 137.835 83.585 ;
        RECT 138.125 83.415 138.295 83.585 ;
        RECT 138.585 83.415 138.755 83.585 ;
        RECT 139.045 83.415 139.215 83.585 ;
        RECT 139.505 83.415 139.675 83.585 ;
        RECT 139.965 83.415 140.135 83.585 ;
        RECT 140.425 83.415 140.595 83.585 ;
        RECT 140.885 83.415 141.055 83.585 ;
        RECT 141.345 83.415 141.515 83.585 ;
        RECT 141.805 83.415 141.975 83.585 ;
        RECT 142.265 83.415 142.435 83.585 ;
        RECT 142.725 83.415 142.895 83.585 ;
        RECT 143.185 83.415 143.355 83.585 ;
        RECT 143.645 83.415 143.815 83.585 ;
        RECT 144.105 83.415 144.275 83.585 ;
        RECT 144.565 83.415 144.735 83.585 ;
        RECT 145.025 83.415 145.195 83.585 ;
        RECT 145.485 83.415 145.655 83.585 ;
        RECT 145.945 83.415 146.115 83.585 ;
        RECT 146.405 83.415 146.575 83.585 ;
        RECT 146.865 83.415 147.035 83.585 ;
        RECT 147.325 83.415 147.495 83.585 ;
        RECT 147.785 83.415 147.955 83.585 ;
        RECT 148.245 83.415 148.415 83.585 ;
        RECT 148.705 83.415 148.875 83.585 ;
        RECT 149.165 83.415 149.335 83.585 ;
        RECT 149.625 83.415 149.795 83.585 ;
        RECT 150.085 83.415 150.255 83.585 ;
        RECT 150.545 83.415 150.715 83.585 ;
        RECT 151.005 83.415 151.175 83.585 ;
        RECT 151.465 83.415 151.635 83.585 ;
        RECT 151.925 83.415 152.095 83.585 ;
        RECT 113.745 82.225 113.915 82.395 ;
        RECT 114.205 81.885 114.375 82.055 ;
        RECT 116.045 82.225 116.215 82.395 ;
        RECT 115.125 81.205 115.295 81.375 ;
        RECT 118.265 82.565 118.435 82.735 ;
        RECT 119.265 82.565 119.435 82.735 ;
        RECT 120.645 82.565 120.815 82.735 ;
        RECT 117.425 81.545 117.595 81.715 ;
        RECT 121.565 82.225 121.735 82.395 ;
        RECT 118.345 81.205 118.515 81.375 ;
        RECT 122.945 82.225 123.115 82.395 ;
        RECT 123.410 82.225 123.580 82.395 ;
        RECT 122.485 81.205 122.655 81.375 ;
        RECT 124.325 81.885 124.495 82.055 ;
        RECT 123.815 81.545 123.985 81.715 ;
        RECT 125.245 82.225 125.415 82.395 ;
        RECT 126.605 82.565 126.775 82.735 ;
        RECT 126.965 82.565 127.135 82.735 ;
        RECT 125.705 81.545 125.875 81.715 ;
        RECT 128.825 82.225 128.995 82.395 ;
        RECT 130.205 82.565 130.375 82.735 ;
        RECT 129.905 82.250 130.075 82.420 ;
        RECT 128.825 81.545 128.995 81.715 ;
        RECT 131.685 81.885 131.855 82.055 ;
        RECT 134.445 82.225 134.615 82.395 ;
        RECT 133.065 81.885 133.235 82.055 ;
        RECT 133.525 81.545 133.695 81.715 ;
        RECT 139.045 82.225 139.215 82.395 ;
        RECT 143.645 82.905 143.815 83.075 ;
        RECT 135.365 81.205 135.535 81.375 ;
        RECT 138.585 81.545 138.755 81.715 ;
        RECT 144.105 82.225 144.275 82.395 ;
        RECT 91.205 80.695 91.375 80.865 ;
        RECT 91.665 80.695 91.835 80.865 ;
        RECT 92.125 80.695 92.295 80.865 ;
        RECT 92.585 80.695 92.755 80.865 ;
        RECT 93.045 80.695 93.215 80.865 ;
        RECT 93.505 80.695 93.675 80.865 ;
        RECT 93.965 80.695 94.135 80.865 ;
        RECT 94.425 80.695 94.595 80.865 ;
        RECT 94.885 80.695 95.055 80.865 ;
        RECT 95.345 80.695 95.515 80.865 ;
        RECT 95.805 80.695 95.975 80.865 ;
        RECT 96.265 80.695 96.435 80.865 ;
        RECT 96.725 80.695 96.895 80.865 ;
        RECT 97.185 80.695 97.355 80.865 ;
        RECT 97.645 80.695 97.815 80.865 ;
        RECT 98.105 80.695 98.275 80.865 ;
        RECT 98.565 80.695 98.735 80.865 ;
        RECT 99.025 80.695 99.195 80.865 ;
        RECT 99.485 80.695 99.655 80.865 ;
        RECT 99.945 80.695 100.115 80.865 ;
        RECT 100.405 80.695 100.575 80.865 ;
        RECT 100.865 80.695 101.035 80.865 ;
        RECT 101.325 80.695 101.495 80.865 ;
        RECT 101.785 80.695 101.955 80.865 ;
        RECT 102.245 80.695 102.415 80.865 ;
        RECT 102.705 80.695 102.875 80.865 ;
        RECT 103.165 80.695 103.335 80.865 ;
        RECT 103.625 80.695 103.795 80.865 ;
        RECT 104.085 80.695 104.255 80.865 ;
        RECT 104.545 80.695 104.715 80.865 ;
        RECT 105.005 80.695 105.175 80.865 ;
        RECT 105.465 80.695 105.635 80.865 ;
        RECT 105.925 80.695 106.095 80.865 ;
        RECT 106.385 80.695 106.555 80.865 ;
        RECT 106.845 80.695 107.015 80.865 ;
        RECT 107.305 80.695 107.475 80.865 ;
        RECT 107.765 80.695 107.935 80.865 ;
        RECT 108.225 80.695 108.395 80.865 ;
        RECT 108.685 80.695 108.855 80.865 ;
        RECT 109.145 80.695 109.315 80.865 ;
        RECT 109.605 80.695 109.775 80.865 ;
        RECT 110.065 80.695 110.235 80.865 ;
        RECT 110.525 80.695 110.695 80.865 ;
        RECT 110.985 80.695 111.155 80.865 ;
        RECT 111.445 80.695 111.615 80.865 ;
        RECT 111.905 80.695 112.075 80.865 ;
        RECT 112.365 80.695 112.535 80.865 ;
        RECT 112.825 80.695 112.995 80.865 ;
        RECT 113.285 80.695 113.455 80.865 ;
        RECT 113.745 80.695 113.915 80.865 ;
        RECT 114.205 80.695 114.375 80.865 ;
        RECT 114.665 80.695 114.835 80.865 ;
        RECT 115.125 80.695 115.295 80.865 ;
        RECT 115.585 80.695 115.755 80.865 ;
        RECT 116.045 80.695 116.215 80.865 ;
        RECT 116.505 80.695 116.675 80.865 ;
        RECT 116.965 80.695 117.135 80.865 ;
        RECT 117.425 80.695 117.595 80.865 ;
        RECT 117.885 80.695 118.055 80.865 ;
        RECT 118.345 80.695 118.515 80.865 ;
        RECT 118.805 80.695 118.975 80.865 ;
        RECT 119.265 80.695 119.435 80.865 ;
        RECT 119.725 80.695 119.895 80.865 ;
        RECT 120.185 80.695 120.355 80.865 ;
        RECT 120.645 80.695 120.815 80.865 ;
        RECT 121.105 80.695 121.275 80.865 ;
        RECT 121.565 80.695 121.735 80.865 ;
        RECT 122.025 80.695 122.195 80.865 ;
        RECT 122.485 80.695 122.655 80.865 ;
        RECT 122.945 80.695 123.115 80.865 ;
        RECT 123.405 80.695 123.575 80.865 ;
        RECT 123.865 80.695 124.035 80.865 ;
        RECT 124.325 80.695 124.495 80.865 ;
        RECT 124.785 80.695 124.955 80.865 ;
        RECT 125.245 80.695 125.415 80.865 ;
        RECT 125.705 80.695 125.875 80.865 ;
        RECT 126.165 80.695 126.335 80.865 ;
        RECT 126.625 80.695 126.795 80.865 ;
        RECT 127.085 80.695 127.255 80.865 ;
        RECT 127.545 80.695 127.715 80.865 ;
        RECT 128.005 80.695 128.175 80.865 ;
        RECT 128.465 80.695 128.635 80.865 ;
        RECT 128.925 80.695 129.095 80.865 ;
        RECT 129.385 80.695 129.555 80.865 ;
        RECT 129.845 80.695 130.015 80.865 ;
        RECT 130.305 80.695 130.475 80.865 ;
        RECT 130.765 80.695 130.935 80.865 ;
        RECT 131.225 80.695 131.395 80.865 ;
        RECT 131.685 80.695 131.855 80.865 ;
        RECT 132.145 80.695 132.315 80.865 ;
        RECT 132.605 80.695 132.775 80.865 ;
        RECT 133.065 80.695 133.235 80.865 ;
        RECT 133.525 80.695 133.695 80.865 ;
        RECT 133.985 80.695 134.155 80.865 ;
        RECT 134.445 80.695 134.615 80.865 ;
        RECT 134.905 80.695 135.075 80.865 ;
        RECT 135.365 80.695 135.535 80.865 ;
        RECT 135.825 80.695 135.995 80.865 ;
        RECT 136.285 80.695 136.455 80.865 ;
        RECT 136.745 80.695 136.915 80.865 ;
        RECT 137.205 80.695 137.375 80.865 ;
        RECT 137.665 80.695 137.835 80.865 ;
        RECT 138.125 80.695 138.295 80.865 ;
        RECT 138.585 80.695 138.755 80.865 ;
        RECT 139.045 80.695 139.215 80.865 ;
        RECT 139.505 80.695 139.675 80.865 ;
        RECT 139.965 80.695 140.135 80.865 ;
        RECT 140.425 80.695 140.595 80.865 ;
        RECT 140.885 80.695 141.055 80.865 ;
        RECT 141.345 80.695 141.515 80.865 ;
        RECT 141.805 80.695 141.975 80.865 ;
        RECT 142.265 80.695 142.435 80.865 ;
        RECT 142.725 80.695 142.895 80.865 ;
        RECT 143.185 80.695 143.355 80.865 ;
        RECT 143.645 80.695 143.815 80.865 ;
        RECT 144.105 80.695 144.275 80.865 ;
        RECT 144.565 80.695 144.735 80.865 ;
        RECT 145.025 80.695 145.195 80.865 ;
        RECT 145.485 80.695 145.655 80.865 ;
        RECT 145.945 80.695 146.115 80.865 ;
        RECT 146.405 80.695 146.575 80.865 ;
        RECT 146.865 80.695 147.035 80.865 ;
        RECT 147.325 80.695 147.495 80.865 ;
        RECT 147.785 80.695 147.955 80.865 ;
        RECT 148.245 80.695 148.415 80.865 ;
        RECT 148.705 80.695 148.875 80.865 ;
        RECT 149.165 80.695 149.335 80.865 ;
        RECT 149.625 80.695 149.795 80.865 ;
        RECT 150.085 80.695 150.255 80.865 ;
        RECT 150.545 80.695 150.715 80.865 ;
        RECT 151.005 80.695 151.175 80.865 ;
        RECT 151.465 80.695 151.635 80.865 ;
        RECT 151.925 80.695 152.095 80.865 ;
        RECT 110.985 79.505 111.155 79.675 ;
        RECT 111.450 79.165 111.620 79.335 ;
        RECT 111.855 79.845 112.025 80.015 ;
        RECT 112.365 78.825 112.535 78.995 ;
        RECT 113.745 79.845 113.915 80.015 ;
        RECT 113.285 79.165 113.455 79.335 ;
        RECT 116.865 79.845 117.035 80.015 ;
        RECT 115.005 78.825 115.175 78.995 ;
        RECT 116.865 79.165 117.035 79.335 ;
        RECT 122.485 80.185 122.655 80.355 ;
        RECT 117.945 79.140 118.115 79.310 ;
        RECT 118.245 78.825 118.415 78.995 ;
        RECT 123.405 79.845 123.575 80.015 ;
        RECT 119.725 78.485 119.895 78.655 ;
        RECT 121.565 78.825 121.735 78.995 ;
        RECT 122.565 78.825 122.735 78.995 ;
        RECT 126.165 79.505 126.335 79.675 ;
        RECT 125.705 79.165 125.875 79.335 ;
        RECT 127.545 79.845 127.715 80.015 ;
        RECT 128.465 80.185 128.635 80.355 ;
        RECT 128.005 79.165 128.175 79.335 ;
        RECT 133.985 80.185 134.155 80.355 ;
        RECT 131.225 79.165 131.395 79.335 ;
        RECT 132.145 78.825 132.315 78.995 ;
        RECT 133.065 79.165 133.235 79.335 ;
        RECT 132.605 78.825 132.775 78.995 ;
        RECT 134.445 79.845 134.615 80.015 ;
        RECT 135.365 79.165 135.535 79.335 ;
        RECT 136.190 79.165 136.360 79.335 ;
        RECT 136.745 79.165 136.915 79.335 ;
        RECT 137.255 79.215 137.425 79.385 ;
        RECT 145.025 80.185 145.195 80.355 ;
        RECT 145.485 79.165 145.655 79.335 ;
        RECT 143.185 78.485 143.355 78.655 ;
        RECT 91.205 77.975 91.375 78.145 ;
        RECT 91.665 77.975 91.835 78.145 ;
        RECT 92.125 77.975 92.295 78.145 ;
        RECT 92.585 77.975 92.755 78.145 ;
        RECT 93.045 77.975 93.215 78.145 ;
        RECT 93.505 77.975 93.675 78.145 ;
        RECT 93.965 77.975 94.135 78.145 ;
        RECT 94.425 77.975 94.595 78.145 ;
        RECT 94.885 77.975 95.055 78.145 ;
        RECT 95.345 77.975 95.515 78.145 ;
        RECT 95.805 77.975 95.975 78.145 ;
        RECT 96.265 77.975 96.435 78.145 ;
        RECT 96.725 77.975 96.895 78.145 ;
        RECT 97.185 77.975 97.355 78.145 ;
        RECT 97.645 77.975 97.815 78.145 ;
        RECT 98.105 77.975 98.275 78.145 ;
        RECT 98.565 77.975 98.735 78.145 ;
        RECT 99.025 77.975 99.195 78.145 ;
        RECT 99.485 77.975 99.655 78.145 ;
        RECT 99.945 77.975 100.115 78.145 ;
        RECT 100.405 77.975 100.575 78.145 ;
        RECT 100.865 77.975 101.035 78.145 ;
        RECT 101.325 77.975 101.495 78.145 ;
        RECT 101.785 77.975 101.955 78.145 ;
        RECT 102.245 77.975 102.415 78.145 ;
        RECT 102.705 77.975 102.875 78.145 ;
        RECT 103.165 77.975 103.335 78.145 ;
        RECT 103.625 77.975 103.795 78.145 ;
        RECT 104.085 77.975 104.255 78.145 ;
        RECT 104.545 77.975 104.715 78.145 ;
        RECT 105.005 77.975 105.175 78.145 ;
        RECT 105.465 77.975 105.635 78.145 ;
        RECT 105.925 77.975 106.095 78.145 ;
        RECT 106.385 77.975 106.555 78.145 ;
        RECT 106.845 77.975 107.015 78.145 ;
        RECT 107.305 77.975 107.475 78.145 ;
        RECT 107.765 77.975 107.935 78.145 ;
        RECT 108.225 77.975 108.395 78.145 ;
        RECT 108.685 77.975 108.855 78.145 ;
        RECT 109.145 77.975 109.315 78.145 ;
        RECT 109.605 77.975 109.775 78.145 ;
        RECT 110.065 77.975 110.235 78.145 ;
        RECT 110.525 77.975 110.695 78.145 ;
        RECT 110.985 77.975 111.155 78.145 ;
        RECT 111.445 77.975 111.615 78.145 ;
        RECT 111.905 77.975 112.075 78.145 ;
        RECT 112.365 77.975 112.535 78.145 ;
        RECT 112.825 77.975 112.995 78.145 ;
        RECT 113.285 77.975 113.455 78.145 ;
        RECT 113.745 77.975 113.915 78.145 ;
        RECT 114.205 77.975 114.375 78.145 ;
        RECT 114.665 77.975 114.835 78.145 ;
        RECT 115.125 77.975 115.295 78.145 ;
        RECT 115.585 77.975 115.755 78.145 ;
        RECT 116.045 77.975 116.215 78.145 ;
        RECT 116.505 77.975 116.675 78.145 ;
        RECT 116.965 77.975 117.135 78.145 ;
        RECT 117.425 77.975 117.595 78.145 ;
        RECT 117.885 77.975 118.055 78.145 ;
        RECT 118.345 77.975 118.515 78.145 ;
        RECT 118.805 77.975 118.975 78.145 ;
        RECT 119.265 77.975 119.435 78.145 ;
        RECT 119.725 77.975 119.895 78.145 ;
        RECT 120.185 77.975 120.355 78.145 ;
        RECT 120.645 77.975 120.815 78.145 ;
        RECT 121.105 77.975 121.275 78.145 ;
        RECT 121.565 77.975 121.735 78.145 ;
        RECT 122.025 77.975 122.195 78.145 ;
        RECT 122.485 77.975 122.655 78.145 ;
        RECT 122.945 77.975 123.115 78.145 ;
        RECT 123.405 77.975 123.575 78.145 ;
        RECT 123.865 77.975 124.035 78.145 ;
        RECT 124.325 77.975 124.495 78.145 ;
        RECT 124.785 77.975 124.955 78.145 ;
        RECT 125.245 77.975 125.415 78.145 ;
        RECT 125.705 77.975 125.875 78.145 ;
        RECT 126.165 77.975 126.335 78.145 ;
        RECT 126.625 77.975 126.795 78.145 ;
        RECT 127.085 77.975 127.255 78.145 ;
        RECT 127.545 77.975 127.715 78.145 ;
        RECT 128.005 77.975 128.175 78.145 ;
        RECT 128.465 77.975 128.635 78.145 ;
        RECT 128.925 77.975 129.095 78.145 ;
        RECT 129.385 77.975 129.555 78.145 ;
        RECT 129.845 77.975 130.015 78.145 ;
        RECT 130.305 77.975 130.475 78.145 ;
        RECT 130.765 77.975 130.935 78.145 ;
        RECT 131.225 77.975 131.395 78.145 ;
        RECT 131.685 77.975 131.855 78.145 ;
        RECT 132.145 77.975 132.315 78.145 ;
        RECT 132.605 77.975 132.775 78.145 ;
        RECT 133.065 77.975 133.235 78.145 ;
        RECT 133.525 77.975 133.695 78.145 ;
        RECT 133.985 77.975 134.155 78.145 ;
        RECT 134.445 77.975 134.615 78.145 ;
        RECT 134.905 77.975 135.075 78.145 ;
        RECT 135.365 77.975 135.535 78.145 ;
        RECT 135.825 77.975 135.995 78.145 ;
        RECT 136.285 77.975 136.455 78.145 ;
        RECT 136.745 77.975 136.915 78.145 ;
        RECT 137.205 77.975 137.375 78.145 ;
        RECT 137.665 77.975 137.835 78.145 ;
        RECT 138.125 77.975 138.295 78.145 ;
        RECT 138.585 77.975 138.755 78.145 ;
        RECT 139.045 77.975 139.215 78.145 ;
        RECT 139.505 77.975 139.675 78.145 ;
        RECT 139.965 77.975 140.135 78.145 ;
        RECT 140.425 77.975 140.595 78.145 ;
        RECT 140.885 77.975 141.055 78.145 ;
        RECT 141.345 77.975 141.515 78.145 ;
        RECT 141.805 77.975 141.975 78.145 ;
        RECT 142.265 77.975 142.435 78.145 ;
        RECT 142.725 77.975 142.895 78.145 ;
        RECT 143.185 77.975 143.355 78.145 ;
        RECT 143.645 77.975 143.815 78.145 ;
        RECT 144.105 77.975 144.275 78.145 ;
        RECT 144.565 77.975 144.735 78.145 ;
        RECT 145.025 77.975 145.195 78.145 ;
        RECT 145.485 77.975 145.655 78.145 ;
        RECT 145.945 77.975 146.115 78.145 ;
        RECT 146.405 77.975 146.575 78.145 ;
        RECT 146.865 77.975 147.035 78.145 ;
        RECT 147.325 77.975 147.495 78.145 ;
        RECT 147.785 77.975 147.955 78.145 ;
        RECT 148.245 77.975 148.415 78.145 ;
        RECT 148.705 77.975 148.875 78.145 ;
        RECT 149.165 77.975 149.335 78.145 ;
        RECT 149.625 77.975 149.795 78.145 ;
        RECT 150.085 77.975 150.255 78.145 ;
        RECT 150.545 77.975 150.715 78.145 ;
        RECT 151.005 77.975 151.175 78.145 ;
        RECT 151.465 77.975 151.635 78.145 ;
        RECT 151.925 77.975 152.095 78.145 ;
        RECT 109.605 76.785 109.775 76.955 ;
        RECT 108.685 75.765 108.855 75.935 ;
        RECT 118.805 77.125 118.975 77.295 ;
        RECT 120.645 77.465 120.815 77.635 ;
        RECT 119.805 77.125 119.975 77.295 ;
        RECT 121.565 77.465 121.735 77.635 ;
        RECT 122.025 76.785 122.195 76.955 ;
        RECT 119.725 75.765 119.895 75.935 ;
        RECT 132.605 76.785 132.775 76.955 ;
        RECT 133.065 76.785 133.235 76.955 ;
        RECT 133.525 76.785 133.695 76.955 ;
        RECT 134.445 77.125 134.615 77.295 ;
        RECT 131.685 75.765 131.855 75.935 ;
        RECT 135.825 76.785 135.995 76.955 ;
        RECT 137.665 76.785 137.835 76.955 ;
        RECT 134.905 75.765 135.075 75.935 ;
        RECT 137.205 75.765 137.375 75.935 ;
        RECT 141.345 75.765 141.515 75.935 ;
        RECT 142.265 76.445 142.435 76.615 ;
        RECT 141.805 75.765 141.975 75.935 ;
        RECT 144.105 76.785 144.275 76.955 ;
        RECT 143.645 76.445 143.815 76.615 ;
        RECT 146.405 76.785 146.575 76.955 ;
        RECT 145.485 75.765 145.655 75.935 ;
        RECT 146.865 75.765 147.035 75.935 ;
        RECT 91.205 75.255 91.375 75.425 ;
        RECT 91.665 75.255 91.835 75.425 ;
        RECT 92.125 75.255 92.295 75.425 ;
        RECT 92.585 75.255 92.755 75.425 ;
        RECT 93.045 75.255 93.215 75.425 ;
        RECT 93.505 75.255 93.675 75.425 ;
        RECT 93.965 75.255 94.135 75.425 ;
        RECT 94.425 75.255 94.595 75.425 ;
        RECT 94.885 75.255 95.055 75.425 ;
        RECT 95.345 75.255 95.515 75.425 ;
        RECT 95.805 75.255 95.975 75.425 ;
        RECT 96.265 75.255 96.435 75.425 ;
        RECT 96.725 75.255 96.895 75.425 ;
        RECT 97.185 75.255 97.355 75.425 ;
        RECT 97.645 75.255 97.815 75.425 ;
        RECT 98.105 75.255 98.275 75.425 ;
        RECT 98.565 75.255 98.735 75.425 ;
        RECT 99.025 75.255 99.195 75.425 ;
        RECT 99.485 75.255 99.655 75.425 ;
        RECT 99.945 75.255 100.115 75.425 ;
        RECT 100.405 75.255 100.575 75.425 ;
        RECT 100.865 75.255 101.035 75.425 ;
        RECT 101.325 75.255 101.495 75.425 ;
        RECT 101.785 75.255 101.955 75.425 ;
        RECT 102.245 75.255 102.415 75.425 ;
        RECT 102.705 75.255 102.875 75.425 ;
        RECT 103.165 75.255 103.335 75.425 ;
        RECT 103.625 75.255 103.795 75.425 ;
        RECT 104.085 75.255 104.255 75.425 ;
        RECT 104.545 75.255 104.715 75.425 ;
        RECT 105.005 75.255 105.175 75.425 ;
        RECT 105.465 75.255 105.635 75.425 ;
        RECT 105.925 75.255 106.095 75.425 ;
        RECT 106.385 75.255 106.555 75.425 ;
        RECT 106.845 75.255 107.015 75.425 ;
        RECT 107.305 75.255 107.475 75.425 ;
        RECT 107.765 75.255 107.935 75.425 ;
        RECT 108.225 75.255 108.395 75.425 ;
        RECT 108.685 75.255 108.855 75.425 ;
        RECT 109.145 75.255 109.315 75.425 ;
        RECT 109.605 75.255 109.775 75.425 ;
        RECT 110.065 75.255 110.235 75.425 ;
        RECT 110.525 75.255 110.695 75.425 ;
        RECT 110.985 75.255 111.155 75.425 ;
        RECT 111.445 75.255 111.615 75.425 ;
        RECT 111.905 75.255 112.075 75.425 ;
        RECT 112.365 75.255 112.535 75.425 ;
        RECT 112.825 75.255 112.995 75.425 ;
        RECT 113.285 75.255 113.455 75.425 ;
        RECT 113.745 75.255 113.915 75.425 ;
        RECT 114.205 75.255 114.375 75.425 ;
        RECT 114.665 75.255 114.835 75.425 ;
        RECT 115.125 75.255 115.295 75.425 ;
        RECT 115.585 75.255 115.755 75.425 ;
        RECT 116.045 75.255 116.215 75.425 ;
        RECT 116.505 75.255 116.675 75.425 ;
        RECT 116.965 75.255 117.135 75.425 ;
        RECT 117.425 75.255 117.595 75.425 ;
        RECT 117.885 75.255 118.055 75.425 ;
        RECT 118.345 75.255 118.515 75.425 ;
        RECT 118.805 75.255 118.975 75.425 ;
        RECT 119.265 75.255 119.435 75.425 ;
        RECT 119.725 75.255 119.895 75.425 ;
        RECT 120.185 75.255 120.355 75.425 ;
        RECT 120.645 75.255 120.815 75.425 ;
        RECT 121.105 75.255 121.275 75.425 ;
        RECT 121.565 75.255 121.735 75.425 ;
        RECT 122.025 75.255 122.195 75.425 ;
        RECT 122.485 75.255 122.655 75.425 ;
        RECT 122.945 75.255 123.115 75.425 ;
        RECT 123.405 75.255 123.575 75.425 ;
        RECT 123.865 75.255 124.035 75.425 ;
        RECT 124.325 75.255 124.495 75.425 ;
        RECT 124.785 75.255 124.955 75.425 ;
        RECT 125.245 75.255 125.415 75.425 ;
        RECT 125.705 75.255 125.875 75.425 ;
        RECT 126.165 75.255 126.335 75.425 ;
        RECT 126.625 75.255 126.795 75.425 ;
        RECT 127.085 75.255 127.255 75.425 ;
        RECT 127.545 75.255 127.715 75.425 ;
        RECT 128.005 75.255 128.175 75.425 ;
        RECT 128.465 75.255 128.635 75.425 ;
        RECT 128.925 75.255 129.095 75.425 ;
        RECT 129.385 75.255 129.555 75.425 ;
        RECT 129.845 75.255 130.015 75.425 ;
        RECT 130.305 75.255 130.475 75.425 ;
        RECT 130.765 75.255 130.935 75.425 ;
        RECT 131.225 75.255 131.395 75.425 ;
        RECT 131.685 75.255 131.855 75.425 ;
        RECT 132.145 75.255 132.315 75.425 ;
        RECT 132.605 75.255 132.775 75.425 ;
        RECT 133.065 75.255 133.235 75.425 ;
        RECT 133.525 75.255 133.695 75.425 ;
        RECT 133.985 75.255 134.155 75.425 ;
        RECT 134.445 75.255 134.615 75.425 ;
        RECT 134.905 75.255 135.075 75.425 ;
        RECT 135.365 75.255 135.535 75.425 ;
        RECT 135.825 75.255 135.995 75.425 ;
        RECT 136.285 75.255 136.455 75.425 ;
        RECT 136.745 75.255 136.915 75.425 ;
        RECT 137.205 75.255 137.375 75.425 ;
        RECT 137.665 75.255 137.835 75.425 ;
        RECT 138.125 75.255 138.295 75.425 ;
        RECT 138.585 75.255 138.755 75.425 ;
        RECT 139.045 75.255 139.215 75.425 ;
        RECT 139.505 75.255 139.675 75.425 ;
        RECT 139.965 75.255 140.135 75.425 ;
        RECT 140.425 75.255 140.595 75.425 ;
        RECT 140.885 75.255 141.055 75.425 ;
        RECT 141.345 75.255 141.515 75.425 ;
        RECT 141.805 75.255 141.975 75.425 ;
        RECT 142.265 75.255 142.435 75.425 ;
        RECT 142.725 75.255 142.895 75.425 ;
        RECT 143.185 75.255 143.355 75.425 ;
        RECT 143.645 75.255 143.815 75.425 ;
        RECT 144.105 75.255 144.275 75.425 ;
        RECT 144.565 75.255 144.735 75.425 ;
        RECT 145.025 75.255 145.195 75.425 ;
        RECT 145.485 75.255 145.655 75.425 ;
        RECT 145.945 75.255 146.115 75.425 ;
        RECT 146.405 75.255 146.575 75.425 ;
        RECT 146.865 75.255 147.035 75.425 ;
        RECT 147.325 75.255 147.495 75.425 ;
        RECT 147.785 75.255 147.955 75.425 ;
        RECT 148.245 75.255 148.415 75.425 ;
        RECT 148.705 75.255 148.875 75.425 ;
        RECT 149.165 75.255 149.335 75.425 ;
        RECT 149.625 75.255 149.795 75.425 ;
        RECT 150.085 75.255 150.255 75.425 ;
        RECT 150.545 75.255 150.715 75.425 ;
        RECT 151.005 75.255 151.175 75.425 ;
        RECT 151.465 75.255 151.635 75.425 ;
        RECT 151.925 75.255 152.095 75.425 ;
        RECT 104.545 74.065 104.715 74.235 ;
        RECT 105.010 73.725 105.180 73.895 ;
        RECT 105.415 74.405 105.585 74.575 ;
        RECT 105.925 73.385 106.095 73.555 ;
        RECT 107.305 74.405 107.475 74.575 ;
        RECT 106.845 73.725 107.015 73.895 ;
        RECT 110.425 74.405 110.595 74.575 ;
        RECT 108.565 73.385 108.735 73.555 ;
        RECT 110.425 73.725 110.595 73.895 ;
        RECT 111.505 73.700 111.675 73.870 ;
        RECT 111.805 73.385 111.975 73.555 ;
        RECT 114.665 73.385 114.835 73.555 ;
        RECT 116.505 74.065 116.675 74.235 ;
        RECT 116.045 73.725 116.215 73.895 ;
        RECT 117.885 73.045 118.055 73.215 ;
        RECT 119.725 74.745 119.895 74.915 ;
        RECT 120.645 73.725 120.815 73.895 ;
        RECT 121.105 74.065 121.275 74.235 ;
        RECT 121.565 73.725 121.735 73.895 ;
        RECT 122.025 73.725 122.195 73.895 ;
        RECT 126.165 74.405 126.335 74.575 ;
        RECT 127.085 73.385 127.255 73.555 ;
        RECT 128.005 73.385 128.175 73.555 ;
        RECT 130.765 74.745 130.935 74.915 ;
        RECT 131.685 73.725 131.855 73.895 ;
        RECT 132.145 73.725 132.315 73.895 ;
        RECT 133.065 73.725 133.235 73.895 ;
        RECT 133.575 73.775 133.745 73.945 ;
        RECT 141.345 74.745 141.515 74.915 ;
        RECT 141.805 73.725 141.975 73.895 ;
        RECT 142.725 73.725 142.895 73.895 ;
        RECT 143.645 73.725 143.815 73.895 ;
        RECT 145.485 73.725 145.655 73.895 ;
        RECT 145.945 73.725 146.115 73.895 ;
        RECT 146.405 73.725 146.575 73.895 ;
        RECT 143.185 73.045 143.355 73.215 ;
        RECT 144.105 73.385 144.275 73.555 ;
        RECT 147.325 73.725 147.495 73.895 ;
        RECT 91.205 72.535 91.375 72.705 ;
        RECT 91.665 72.535 91.835 72.705 ;
        RECT 92.125 72.535 92.295 72.705 ;
        RECT 92.585 72.535 92.755 72.705 ;
        RECT 93.045 72.535 93.215 72.705 ;
        RECT 93.505 72.535 93.675 72.705 ;
        RECT 93.965 72.535 94.135 72.705 ;
        RECT 94.425 72.535 94.595 72.705 ;
        RECT 94.885 72.535 95.055 72.705 ;
        RECT 95.345 72.535 95.515 72.705 ;
        RECT 95.805 72.535 95.975 72.705 ;
        RECT 96.265 72.535 96.435 72.705 ;
        RECT 96.725 72.535 96.895 72.705 ;
        RECT 97.185 72.535 97.355 72.705 ;
        RECT 97.645 72.535 97.815 72.705 ;
        RECT 98.105 72.535 98.275 72.705 ;
        RECT 98.565 72.535 98.735 72.705 ;
        RECT 99.025 72.535 99.195 72.705 ;
        RECT 99.485 72.535 99.655 72.705 ;
        RECT 99.945 72.535 100.115 72.705 ;
        RECT 100.405 72.535 100.575 72.705 ;
        RECT 100.865 72.535 101.035 72.705 ;
        RECT 101.325 72.535 101.495 72.705 ;
        RECT 101.785 72.535 101.955 72.705 ;
        RECT 102.245 72.535 102.415 72.705 ;
        RECT 102.705 72.535 102.875 72.705 ;
        RECT 103.165 72.535 103.335 72.705 ;
        RECT 103.625 72.535 103.795 72.705 ;
        RECT 104.085 72.535 104.255 72.705 ;
        RECT 104.545 72.535 104.715 72.705 ;
        RECT 105.005 72.535 105.175 72.705 ;
        RECT 105.465 72.535 105.635 72.705 ;
        RECT 105.925 72.535 106.095 72.705 ;
        RECT 106.385 72.535 106.555 72.705 ;
        RECT 106.845 72.535 107.015 72.705 ;
        RECT 107.305 72.535 107.475 72.705 ;
        RECT 107.765 72.535 107.935 72.705 ;
        RECT 108.225 72.535 108.395 72.705 ;
        RECT 108.685 72.535 108.855 72.705 ;
        RECT 109.145 72.535 109.315 72.705 ;
        RECT 109.605 72.535 109.775 72.705 ;
        RECT 110.065 72.535 110.235 72.705 ;
        RECT 110.525 72.535 110.695 72.705 ;
        RECT 110.985 72.535 111.155 72.705 ;
        RECT 111.445 72.535 111.615 72.705 ;
        RECT 111.905 72.535 112.075 72.705 ;
        RECT 112.365 72.535 112.535 72.705 ;
        RECT 112.825 72.535 112.995 72.705 ;
        RECT 113.285 72.535 113.455 72.705 ;
        RECT 113.745 72.535 113.915 72.705 ;
        RECT 114.205 72.535 114.375 72.705 ;
        RECT 114.665 72.535 114.835 72.705 ;
        RECT 115.125 72.535 115.295 72.705 ;
        RECT 115.585 72.535 115.755 72.705 ;
        RECT 116.045 72.535 116.215 72.705 ;
        RECT 116.505 72.535 116.675 72.705 ;
        RECT 116.965 72.535 117.135 72.705 ;
        RECT 117.425 72.535 117.595 72.705 ;
        RECT 117.885 72.535 118.055 72.705 ;
        RECT 118.345 72.535 118.515 72.705 ;
        RECT 118.805 72.535 118.975 72.705 ;
        RECT 119.265 72.535 119.435 72.705 ;
        RECT 119.725 72.535 119.895 72.705 ;
        RECT 120.185 72.535 120.355 72.705 ;
        RECT 120.645 72.535 120.815 72.705 ;
        RECT 121.105 72.535 121.275 72.705 ;
        RECT 121.565 72.535 121.735 72.705 ;
        RECT 122.025 72.535 122.195 72.705 ;
        RECT 122.485 72.535 122.655 72.705 ;
        RECT 122.945 72.535 123.115 72.705 ;
        RECT 123.405 72.535 123.575 72.705 ;
        RECT 123.865 72.535 124.035 72.705 ;
        RECT 124.325 72.535 124.495 72.705 ;
        RECT 124.785 72.535 124.955 72.705 ;
        RECT 125.245 72.535 125.415 72.705 ;
        RECT 125.705 72.535 125.875 72.705 ;
        RECT 126.165 72.535 126.335 72.705 ;
        RECT 126.625 72.535 126.795 72.705 ;
        RECT 127.085 72.535 127.255 72.705 ;
        RECT 127.545 72.535 127.715 72.705 ;
        RECT 128.005 72.535 128.175 72.705 ;
        RECT 128.465 72.535 128.635 72.705 ;
        RECT 128.925 72.535 129.095 72.705 ;
        RECT 129.385 72.535 129.555 72.705 ;
        RECT 129.845 72.535 130.015 72.705 ;
        RECT 130.305 72.535 130.475 72.705 ;
        RECT 130.765 72.535 130.935 72.705 ;
        RECT 131.225 72.535 131.395 72.705 ;
        RECT 131.685 72.535 131.855 72.705 ;
        RECT 132.145 72.535 132.315 72.705 ;
        RECT 132.605 72.535 132.775 72.705 ;
        RECT 133.065 72.535 133.235 72.705 ;
        RECT 133.525 72.535 133.695 72.705 ;
        RECT 133.985 72.535 134.155 72.705 ;
        RECT 134.445 72.535 134.615 72.705 ;
        RECT 134.905 72.535 135.075 72.705 ;
        RECT 135.365 72.535 135.535 72.705 ;
        RECT 135.825 72.535 135.995 72.705 ;
        RECT 136.285 72.535 136.455 72.705 ;
        RECT 136.745 72.535 136.915 72.705 ;
        RECT 137.205 72.535 137.375 72.705 ;
        RECT 137.665 72.535 137.835 72.705 ;
        RECT 138.125 72.535 138.295 72.705 ;
        RECT 138.585 72.535 138.755 72.705 ;
        RECT 139.045 72.535 139.215 72.705 ;
        RECT 139.505 72.535 139.675 72.705 ;
        RECT 139.965 72.535 140.135 72.705 ;
        RECT 140.425 72.535 140.595 72.705 ;
        RECT 140.885 72.535 141.055 72.705 ;
        RECT 141.345 72.535 141.515 72.705 ;
        RECT 141.805 72.535 141.975 72.705 ;
        RECT 142.265 72.535 142.435 72.705 ;
        RECT 142.725 72.535 142.895 72.705 ;
        RECT 143.185 72.535 143.355 72.705 ;
        RECT 143.645 72.535 143.815 72.705 ;
        RECT 144.105 72.535 144.275 72.705 ;
        RECT 144.565 72.535 144.735 72.705 ;
        RECT 145.025 72.535 145.195 72.705 ;
        RECT 145.485 72.535 145.655 72.705 ;
        RECT 145.945 72.535 146.115 72.705 ;
        RECT 146.405 72.535 146.575 72.705 ;
        RECT 146.865 72.535 147.035 72.705 ;
        RECT 147.325 72.535 147.495 72.705 ;
        RECT 147.785 72.535 147.955 72.705 ;
        RECT 148.245 72.535 148.415 72.705 ;
        RECT 148.705 72.535 148.875 72.705 ;
        RECT 149.165 72.535 149.335 72.705 ;
        RECT 149.625 72.535 149.795 72.705 ;
        RECT 150.085 72.535 150.255 72.705 ;
        RECT 150.545 72.535 150.715 72.705 ;
        RECT 151.005 72.535 151.175 72.705 ;
        RECT 151.465 72.535 151.635 72.705 ;
        RECT 151.925 72.535 152.095 72.705 ;
        RECT 23.500 71.940 23.760 72.200 ;
        RECT 32.960 71.970 33.340 72.280 ;
        RECT 21.890 69.410 22.060 70.290 ;
        RECT 22.330 69.410 22.500 70.290 ;
        RECT 21.890 67.740 22.060 68.620 ;
        RECT 22.330 67.740 22.500 68.620 ;
        RECT 20.125 67.030 20.330 67.230 ;
        RECT 24.310 69.690 24.480 70.570 ;
        RECT 24.310 67.740 24.480 68.620 ;
        RECT 24.750 69.690 24.920 70.570 ;
        RECT 24.750 67.740 24.920 68.620 ;
        RECT 25.190 69.690 25.360 70.570 ;
        RECT 25.190 67.740 25.360 68.620 ;
        RECT 21.900 65.450 22.070 66.330 ;
        RECT 26.180 69.000 26.350 69.880 ;
        RECT 26.620 69.000 26.790 69.880 ;
        RECT 27.570 69.705 27.905 70.030 ;
        RECT 26.180 67.330 26.350 68.210 ;
        RECT 26.620 67.330 26.790 68.210 ;
        RECT 27.470 67.450 27.770 67.740 ;
        RECT 22.340 65.450 22.510 66.330 ;
        RECT 21.900 63.780 22.070 64.660 ;
        RECT 22.340 63.780 22.510 64.660 ;
        RECT 23.540 65.410 23.710 66.290 ;
        RECT 19.080 63.390 19.420 63.660 ;
        RECT 23.540 63.460 23.710 64.340 ;
        RECT 21.495 61.895 21.760 62.115 ;
        RECT 23.980 65.410 24.150 66.290 ;
        RECT 23.980 63.460 24.150 64.340 ;
        RECT 24.420 65.410 24.590 66.290 ;
        RECT 24.420 63.460 24.590 64.340 ;
        RECT 25.070 65.410 25.240 66.290 ;
        RECT 25.070 63.460 25.240 64.340 ;
        RECT 25.510 65.410 25.680 66.290 ;
        RECT 25.510 63.460 25.680 64.340 ;
        RECT 25.950 65.410 26.120 66.290 ;
        RECT 25.950 63.460 26.120 64.340 ;
        RECT 26.560 65.410 26.730 66.290 ;
        RECT 27.000 65.410 27.170 66.290 ;
        RECT 29.640 69.690 29.810 70.570 ;
        RECT 29.640 67.740 29.810 68.620 ;
        RECT 30.080 69.690 30.250 70.570 ;
        RECT 30.080 67.740 30.250 68.620 ;
        RECT 30.520 69.690 30.690 70.570 ;
        RECT 31.140 69.240 31.310 69.415 ;
        RECT 31.750 69.000 31.920 69.880 ;
        RECT 34.380 70.220 34.550 70.395 ;
        RECT 32.190 69.000 32.360 69.880 ;
        RECT 30.520 67.740 30.690 68.620 ;
        RECT 31.750 67.330 31.920 68.210 ;
        RECT 32.190 67.330 32.360 68.210 ;
        RECT 32.800 69.000 32.970 69.880 ;
        RECT 33.240 69.000 33.410 69.880 ;
        RECT 109.145 72.025 109.315 72.195 ;
        RECT 108.685 71.345 108.855 71.515 ;
        RECT 115.125 71.345 115.295 71.515 ;
        RECT 117.425 72.025 117.595 72.195 ;
        RECT 116.045 71.345 116.215 71.515 ;
        RECT 116.505 71.345 116.675 71.515 ;
        RECT 115.125 70.325 115.295 70.495 ;
        RECT 117.885 70.665 118.055 70.835 ;
        RECT 119.725 71.685 119.895 71.855 ;
        RECT 122.025 71.005 122.195 71.175 ;
        RECT 125.705 72.025 125.875 72.195 ;
        RECT 124.785 71.345 124.955 71.515 ;
        RECT 125.245 71.345 125.415 71.515 ;
        RECT 126.165 71.345 126.335 71.515 ;
        RECT 126.625 71.345 126.795 71.515 ;
        RECT 127.545 71.685 127.715 71.855 ;
        RECT 128.005 71.345 128.175 71.515 ;
        RECT 133.525 71.685 133.695 71.855 ;
        RECT 126.625 70.325 126.795 70.495 ;
        RECT 134.445 71.345 134.615 71.515 ;
        RECT 134.905 70.665 135.075 70.835 ;
        RECT 135.365 71.345 135.535 71.515 ;
        RECT 135.825 71.345 135.995 71.515 ;
        RECT 139.045 72.025 139.215 72.195 ;
        RECT 137.665 71.345 137.835 71.515 ;
        RECT 139.505 71.345 139.675 71.515 ;
        RECT 137.205 70.325 137.375 70.495 ;
        RECT 141.345 70.665 141.515 70.835 ;
        RECT 142.265 70.665 142.435 70.835 ;
        RECT 143.185 70.665 143.355 70.835 ;
        RECT 145.025 72.025 145.195 72.195 ;
        RECT 145.945 70.665 146.115 70.835 ;
        RECT 145.025 70.325 145.195 70.495 ;
        RECT 149.165 71.345 149.335 71.515 ;
        RECT 150.545 71.005 150.715 71.175 ;
        RECT 91.205 69.815 91.375 69.985 ;
        RECT 91.665 69.815 91.835 69.985 ;
        RECT 92.125 69.815 92.295 69.985 ;
        RECT 92.585 69.815 92.755 69.985 ;
        RECT 93.045 69.815 93.215 69.985 ;
        RECT 93.505 69.815 93.675 69.985 ;
        RECT 93.965 69.815 94.135 69.985 ;
        RECT 94.425 69.815 94.595 69.985 ;
        RECT 94.885 69.815 95.055 69.985 ;
        RECT 95.345 69.815 95.515 69.985 ;
        RECT 95.805 69.815 95.975 69.985 ;
        RECT 96.265 69.815 96.435 69.985 ;
        RECT 96.725 69.815 96.895 69.985 ;
        RECT 97.185 69.815 97.355 69.985 ;
        RECT 97.645 69.815 97.815 69.985 ;
        RECT 98.105 69.815 98.275 69.985 ;
        RECT 98.565 69.815 98.735 69.985 ;
        RECT 99.025 69.815 99.195 69.985 ;
        RECT 99.485 69.815 99.655 69.985 ;
        RECT 99.945 69.815 100.115 69.985 ;
        RECT 100.405 69.815 100.575 69.985 ;
        RECT 100.865 69.815 101.035 69.985 ;
        RECT 101.325 69.815 101.495 69.985 ;
        RECT 101.785 69.815 101.955 69.985 ;
        RECT 102.245 69.815 102.415 69.985 ;
        RECT 102.705 69.815 102.875 69.985 ;
        RECT 103.165 69.815 103.335 69.985 ;
        RECT 103.625 69.815 103.795 69.985 ;
        RECT 104.085 69.815 104.255 69.985 ;
        RECT 104.545 69.815 104.715 69.985 ;
        RECT 105.005 69.815 105.175 69.985 ;
        RECT 105.465 69.815 105.635 69.985 ;
        RECT 105.925 69.815 106.095 69.985 ;
        RECT 106.385 69.815 106.555 69.985 ;
        RECT 106.845 69.815 107.015 69.985 ;
        RECT 107.305 69.815 107.475 69.985 ;
        RECT 107.765 69.815 107.935 69.985 ;
        RECT 108.225 69.815 108.395 69.985 ;
        RECT 108.685 69.815 108.855 69.985 ;
        RECT 109.145 69.815 109.315 69.985 ;
        RECT 109.605 69.815 109.775 69.985 ;
        RECT 110.065 69.815 110.235 69.985 ;
        RECT 110.525 69.815 110.695 69.985 ;
        RECT 110.985 69.815 111.155 69.985 ;
        RECT 111.445 69.815 111.615 69.985 ;
        RECT 111.905 69.815 112.075 69.985 ;
        RECT 112.365 69.815 112.535 69.985 ;
        RECT 112.825 69.815 112.995 69.985 ;
        RECT 113.285 69.815 113.455 69.985 ;
        RECT 113.745 69.815 113.915 69.985 ;
        RECT 114.205 69.815 114.375 69.985 ;
        RECT 114.665 69.815 114.835 69.985 ;
        RECT 115.125 69.815 115.295 69.985 ;
        RECT 115.585 69.815 115.755 69.985 ;
        RECT 116.045 69.815 116.215 69.985 ;
        RECT 116.505 69.815 116.675 69.985 ;
        RECT 116.965 69.815 117.135 69.985 ;
        RECT 117.425 69.815 117.595 69.985 ;
        RECT 117.885 69.815 118.055 69.985 ;
        RECT 118.345 69.815 118.515 69.985 ;
        RECT 118.805 69.815 118.975 69.985 ;
        RECT 119.265 69.815 119.435 69.985 ;
        RECT 119.725 69.815 119.895 69.985 ;
        RECT 120.185 69.815 120.355 69.985 ;
        RECT 120.645 69.815 120.815 69.985 ;
        RECT 121.105 69.815 121.275 69.985 ;
        RECT 121.565 69.815 121.735 69.985 ;
        RECT 122.025 69.815 122.195 69.985 ;
        RECT 122.485 69.815 122.655 69.985 ;
        RECT 122.945 69.815 123.115 69.985 ;
        RECT 123.405 69.815 123.575 69.985 ;
        RECT 123.865 69.815 124.035 69.985 ;
        RECT 124.325 69.815 124.495 69.985 ;
        RECT 124.785 69.815 124.955 69.985 ;
        RECT 125.245 69.815 125.415 69.985 ;
        RECT 125.705 69.815 125.875 69.985 ;
        RECT 126.165 69.815 126.335 69.985 ;
        RECT 126.625 69.815 126.795 69.985 ;
        RECT 127.085 69.815 127.255 69.985 ;
        RECT 127.545 69.815 127.715 69.985 ;
        RECT 128.005 69.815 128.175 69.985 ;
        RECT 128.465 69.815 128.635 69.985 ;
        RECT 128.925 69.815 129.095 69.985 ;
        RECT 129.385 69.815 129.555 69.985 ;
        RECT 129.845 69.815 130.015 69.985 ;
        RECT 130.305 69.815 130.475 69.985 ;
        RECT 130.765 69.815 130.935 69.985 ;
        RECT 131.225 69.815 131.395 69.985 ;
        RECT 131.685 69.815 131.855 69.985 ;
        RECT 132.145 69.815 132.315 69.985 ;
        RECT 132.605 69.815 132.775 69.985 ;
        RECT 133.065 69.815 133.235 69.985 ;
        RECT 133.525 69.815 133.695 69.985 ;
        RECT 133.985 69.815 134.155 69.985 ;
        RECT 134.445 69.815 134.615 69.985 ;
        RECT 134.905 69.815 135.075 69.985 ;
        RECT 135.365 69.815 135.535 69.985 ;
        RECT 135.825 69.815 135.995 69.985 ;
        RECT 136.285 69.815 136.455 69.985 ;
        RECT 136.745 69.815 136.915 69.985 ;
        RECT 137.205 69.815 137.375 69.985 ;
        RECT 137.665 69.815 137.835 69.985 ;
        RECT 138.125 69.815 138.295 69.985 ;
        RECT 138.585 69.815 138.755 69.985 ;
        RECT 139.045 69.815 139.215 69.985 ;
        RECT 139.505 69.815 139.675 69.985 ;
        RECT 139.965 69.815 140.135 69.985 ;
        RECT 140.425 69.815 140.595 69.985 ;
        RECT 140.885 69.815 141.055 69.985 ;
        RECT 141.345 69.815 141.515 69.985 ;
        RECT 141.805 69.815 141.975 69.985 ;
        RECT 142.265 69.815 142.435 69.985 ;
        RECT 142.725 69.815 142.895 69.985 ;
        RECT 143.185 69.815 143.355 69.985 ;
        RECT 143.645 69.815 143.815 69.985 ;
        RECT 144.105 69.815 144.275 69.985 ;
        RECT 144.565 69.815 144.735 69.985 ;
        RECT 145.025 69.815 145.195 69.985 ;
        RECT 145.485 69.815 145.655 69.985 ;
        RECT 145.945 69.815 146.115 69.985 ;
        RECT 146.405 69.815 146.575 69.985 ;
        RECT 146.865 69.815 147.035 69.985 ;
        RECT 147.325 69.815 147.495 69.985 ;
        RECT 147.785 69.815 147.955 69.985 ;
        RECT 148.245 69.815 148.415 69.985 ;
        RECT 148.705 69.815 148.875 69.985 ;
        RECT 149.165 69.815 149.335 69.985 ;
        RECT 149.625 69.815 149.795 69.985 ;
        RECT 150.085 69.815 150.255 69.985 ;
        RECT 150.545 69.815 150.715 69.985 ;
        RECT 151.005 69.815 151.175 69.985 ;
        RECT 151.465 69.815 151.635 69.985 ;
        RECT 151.925 69.815 152.095 69.985 ;
        RECT 32.800 67.330 32.970 68.210 ;
        RECT 31.745 66.705 31.915 66.875 ;
        RECT 28.870 65.410 29.040 66.290 ;
        RECT 26.560 63.740 26.730 64.620 ;
        RECT 27.000 63.740 27.170 64.620 ;
        RECT 25.035 59.445 25.320 59.670 ;
        RECT 6.110 56.755 6.300 58.740 ;
        RECT 27.730 63.340 28.065 63.665 ;
        RECT 28.870 63.460 29.040 64.340 ;
        RECT 29.310 65.410 29.480 66.290 ;
        RECT 29.310 63.460 29.480 64.340 ;
        RECT 29.750 65.410 29.920 66.290 ;
        RECT 29.750 63.460 29.920 64.340 ;
        RECT 30.400 65.410 30.570 66.290 ;
        RECT 30.400 63.460 30.570 64.340 ;
        RECT 28.780 59.195 29.190 59.545 ;
        RECT 30.840 65.410 31.010 66.290 ;
        RECT 30.840 63.460 31.010 64.340 ;
        RECT 31.280 65.410 31.450 66.290 ;
        RECT 33.240 67.330 33.410 68.210 ;
        RECT 33.965 66.710 34.150 66.910 ;
        RECT 32.095 65.350 32.265 66.230 ;
        RECT 32.535 65.350 32.705 66.230 ;
        RECT 31.280 63.460 31.450 64.340 ;
        RECT 31.175 62.425 31.350 62.600 ;
        RECT 32.095 63.680 32.265 64.560 ;
        RECT 32.535 63.680 32.705 64.560 ;
        RECT 33.145 65.350 33.315 66.230 ;
        RECT 33.585 65.350 33.755 66.230 ;
        RECT 102.245 68.285 102.415 68.455 ;
        RECT 101.325 67.605 101.495 67.775 ;
        RECT 110.985 68.625 111.155 68.795 ;
        RECT 111.450 68.285 111.620 68.455 ;
        RECT 111.855 68.965 112.025 69.135 ;
        RECT 112.365 68.625 112.535 68.795 ;
        RECT 113.745 68.965 113.915 69.135 ;
        RECT 113.285 68.285 113.455 68.455 ;
        RECT 116.865 68.965 117.035 69.135 ;
        RECT 115.005 67.945 115.175 68.115 ;
        RECT 116.865 68.285 117.035 68.455 ;
        RECT 119.725 68.625 119.895 68.795 ;
        RECT 120.645 69.305 120.815 69.475 ;
        RECT 117.945 68.260 118.115 68.430 ;
        RECT 118.245 67.945 118.415 68.115 ;
        RECT 121.565 68.285 121.735 68.455 ;
        RECT 122.485 68.285 122.655 68.455 ;
        RECT 132.145 68.625 132.315 68.795 ;
        RECT 134.445 69.305 134.615 69.475 ;
        RECT 133.985 68.965 134.155 69.135 ;
        RECT 135.365 69.305 135.535 69.475 ;
        RECT 138.125 69.305 138.295 69.475 ;
        RECT 134.905 68.285 135.075 68.455 ;
        RECT 139.965 69.305 140.135 69.475 ;
        RECT 137.665 68.285 137.835 68.455 ;
        RECT 137.205 67.605 137.375 67.775 ;
        RECT 145.945 69.305 146.115 69.475 ;
        RECT 142.725 68.285 142.895 68.455 ;
        RECT 143.190 68.285 143.360 68.455 ;
        RECT 144.105 67.945 144.275 68.115 ;
        RECT 145.050 68.285 145.220 68.455 ;
        RECT 144.565 67.945 144.735 68.115 ;
        RECT 147.325 69.305 147.495 69.475 ;
        RECT 146.405 68.625 146.575 68.795 ;
        RECT 148.705 68.285 148.875 68.455 ;
        RECT 91.205 67.095 91.375 67.265 ;
        RECT 91.665 67.095 91.835 67.265 ;
        RECT 92.125 67.095 92.295 67.265 ;
        RECT 92.585 67.095 92.755 67.265 ;
        RECT 93.045 67.095 93.215 67.265 ;
        RECT 93.505 67.095 93.675 67.265 ;
        RECT 93.965 67.095 94.135 67.265 ;
        RECT 94.425 67.095 94.595 67.265 ;
        RECT 94.885 67.095 95.055 67.265 ;
        RECT 95.345 67.095 95.515 67.265 ;
        RECT 95.805 67.095 95.975 67.265 ;
        RECT 96.265 67.095 96.435 67.265 ;
        RECT 96.725 67.095 96.895 67.265 ;
        RECT 97.185 67.095 97.355 67.265 ;
        RECT 97.645 67.095 97.815 67.265 ;
        RECT 98.105 67.095 98.275 67.265 ;
        RECT 98.565 67.095 98.735 67.265 ;
        RECT 99.025 67.095 99.195 67.265 ;
        RECT 99.485 67.095 99.655 67.265 ;
        RECT 99.945 67.095 100.115 67.265 ;
        RECT 100.405 67.095 100.575 67.265 ;
        RECT 100.865 67.095 101.035 67.265 ;
        RECT 101.325 67.095 101.495 67.265 ;
        RECT 101.785 67.095 101.955 67.265 ;
        RECT 102.245 67.095 102.415 67.265 ;
        RECT 102.705 67.095 102.875 67.265 ;
        RECT 103.165 67.095 103.335 67.265 ;
        RECT 103.625 67.095 103.795 67.265 ;
        RECT 104.085 67.095 104.255 67.265 ;
        RECT 104.545 67.095 104.715 67.265 ;
        RECT 105.005 67.095 105.175 67.265 ;
        RECT 105.465 67.095 105.635 67.265 ;
        RECT 105.925 67.095 106.095 67.265 ;
        RECT 106.385 67.095 106.555 67.265 ;
        RECT 106.845 67.095 107.015 67.265 ;
        RECT 107.305 67.095 107.475 67.265 ;
        RECT 107.765 67.095 107.935 67.265 ;
        RECT 108.225 67.095 108.395 67.265 ;
        RECT 108.685 67.095 108.855 67.265 ;
        RECT 109.145 67.095 109.315 67.265 ;
        RECT 109.605 67.095 109.775 67.265 ;
        RECT 110.065 67.095 110.235 67.265 ;
        RECT 110.525 67.095 110.695 67.265 ;
        RECT 110.985 67.095 111.155 67.265 ;
        RECT 111.445 67.095 111.615 67.265 ;
        RECT 111.905 67.095 112.075 67.265 ;
        RECT 112.365 67.095 112.535 67.265 ;
        RECT 112.825 67.095 112.995 67.265 ;
        RECT 113.285 67.095 113.455 67.265 ;
        RECT 113.745 67.095 113.915 67.265 ;
        RECT 114.205 67.095 114.375 67.265 ;
        RECT 114.665 67.095 114.835 67.265 ;
        RECT 115.125 67.095 115.295 67.265 ;
        RECT 115.585 67.095 115.755 67.265 ;
        RECT 116.045 67.095 116.215 67.265 ;
        RECT 116.505 67.095 116.675 67.265 ;
        RECT 116.965 67.095 117.135 67.265 ;
        RECT 117.425 67.095 117.595 67.265 ;
        RECT 117.885 67.095 118.055 67.265 ;
        RECT 118.345 67.095 118.515 67.265 ;
        RECT 118.805 67.095 118.975 67.265 ;
        RECT 119.265 67.095 119.435 67.265 ;
        RECT 119.725 67.095 119.895 67.265 ;
        RECT 120.185 67.095 120.355 67.265 ;
        RECT 120.645 67.095 120.815 67.265 ;
        RECT 121.105 67.095 121.275 67.265 ;
        RECT 121.565 67.095 121.735 67.265 ;
        RECT 122.025 67.095 122.195 67.265 ;
        RECT 122.485 67.095 122.655 67.265 ;
        RECT 122.945 67.095 123.115 67.265 ;
        RECT 123.405 67.095 123.575 67.265 ;
        RECT 123.865 67.095 124.035 67.265 ;
        RECT 124.325 67.095 124.495 67.265 ;
        RECT 124.785 67.095 124.955 67.265 ;
        RECT 125.245 67.095 125.415 67.265 ;
        RECT 125.705 67.095 125.875 67.265 ;
        RECT 126.165 67.095 126.335 67.265 ;
        RECT 126.625 67.095 126.795 67.265 ;
        RECT 127.085 67.095 127.255 67.265 ;
        RECT 127.545 67.095 127.715 67.265 ;
        RECT 128.005 67.095 128.175 67.265 ;
        RECT 128.465 67.095 128.635 67.265 ;
        RECT 128.925 67.095 129.095 67.265 ;
        RECT 129.385 67.095 129.555 67.265 ;
        RECT 129.845 67.095 130.015 67.265 ;
        RECT 130.305 67.095 130.475 67.265 ;
        RECT 130.765 67.095 130.935 67.265 ;
        RECT 131.225 67.095 131.395 67.265 ;
        RECT 131.685 67.095 131.855 67.265 ;
        RECT 132.145 67.095 132.315 67.265 ;
        RECT 132.605 67.095 132.775 67.265 ;
        RECT 133.065 67.095 133.235 67.265 ;
        RECT 133.525 67.095 133.695 67.265 ;
        RECT 133.985 67.095 134.155 67.265 ;
        RECT 134.445 67.095 134.615 67.265 ;
        RECT 134.905 67.095 135.075 67.265 ;
        RECT 135.365 67.095 135.535 67.265 ;
        RECT 135.825 67.095 135.995 67.265 ;
        RECT 136.285 67.095 136.455 67.265 ;
        RECT 136.745 67.095 136.915 67.265 ;
        RECT 137.205 67.095 137.375 67.265 ;
        RECT 137.665 67.095 137.835 67.265 ;
        RECT 138.125 67.095 138.295 67.265 ;
        RECT 138.585 67.095 138.755 67.265 ;
        RECT 139.045 67.095 139.215 67.265 ;
        RECT 139.505 67.095 139.675 67.265 ;
        RECT 139.965 67.095 140.135 67.265 ;
        RECT 140.425 67.095 140.595 67.265 ;
        RECT 140.885 67.095 141.055 67.265 ;
        RECT 141.345 67.095 141.515 67.265 ;
        RECT 141.805 67.095 141.975 67.265 ;
        RECT 142.265 67.095 142.435 67.265 ;
        RECT 142.725 67.095 142.895 67.265 ;
        RECT 143.185 67.095 143.355 67.265 ;
        RECT 143.645 67.095 143.815 67.265 ;
        RECT 144.105 67.095 144.275 67.265 ;
        RECT 144.565 67.095 144.735 67.265 ;
        RECT 145.025 67.095 145.195 67.265 ;
        RECT 145.485 67.095 145.655 67.265 ;
        RECT 145.945 67.095 146.115 67.265 ;
        RECT 146.405 67.095 146.575 67.265 ;
        RECT 146.865 67.095 147.035 67.265 ;
        RECT 147.325 67.095 147.495 67.265 ;
        RECT 147.785 67.095 147.955 67.265 ;
        RECT 148.245 67.095 148.415 67.265 ;
        RECT 148.705 67.095 148.875 67.265 ;
        RECT 149.165 67.095 149.335 67.265 ;
        RECT 149.625 67.095 149.795 67.265 ;
        RECT 150.085 67.095 150.255 67.265 ;
        RECT 150.545 67.095 150.715 67.265 ;
        RECT 151.005 67.095 151.175 67.265 ;
        RECT 151.465 67.095 151.635 67.265 ;
        RECT 151.925 67.095 152.095 67.265 ;
        RECT 35.225 65.665 35.495 65.925 ;
        RECT 34.540 64.690 34.850 64.970 ;
        RECT 33.145 63.680 33.315 64.560 ;
        RECT 33.585 63.680 33.755 64.560 ;
        RECT 98.565 65.565 98.735 65.735 ;
        RECT 99.030 65.905 99.200 66.075 ;
        RECT 99.945 66.245 100.115 66.415 ;
        RECT 99.435 65.225 99.605 65.395 ;
        RECT 100.865 65.905 101.035 66.075 ;
        RECT 102.225 66.245 102.395 66.415 ;
        RECT 102.585 66.245 102.755 66.415 ;
        RECT 101.325 65.225 101.495 65.395 ;
        RECT 104.445 65.905 104.615 66.075 ;
        RECT 105.825 66.245 105.995 66.415 ;
        RECT 105.525 65.930 105.695 66.100 ;
        RECT 104.445 65.225 104.615 65.395 ;
        RECT 108.685 66.245 108.855 66.415 ;
        RECT 109.145 65.905 109.315 66.075 ;
        RECT 115.585 66.245 115.755 66.415 ;
        RECT 107.305 64.885 107.475 65.055 ;
        RECT 115.125 65.905 115.295 66.075 ;
        RECT 122.945 65.905 123.115 66.075 ;
        RECT 124.325 65.905 124.495 66.075 ;
        RECT 122.485 64.885 122.655 65.055 ;
        RECT 124.790 65.905 124.960 66.075 ;
        RECT 125.705 65.565 125.875 65.735 ;
        RECT 125.195 65.225 125.365 65.395 ;
        RECT 126.625 65.905 126.795 66.075 ;
        RECT 127.985 66.245 128.155 66.415 ;
        RECT 128.345 66.245 128.515 66.415 ;
        RECT 127.085 65.225 127.255 65.395 ;
        RECT 130.205 65.905 130.375 66.075 ;
        RECT 131.585 66.245 131.755 66.415 ;
        RECT 131.285 65.930 131.455 66.100 ;
        RECT 130.205 65.225 130.375 65.395 ;
        RECT 135.365 66.245 135.535 66.415 ;
        RECT 134.445 65.905 134.615 66.075 ;
        RECT 133.065 65.565 133.235 65.735 ;
        RECT 135.365 65.565 135.535 65.735 ;
        RECT 139.505 65.905 139.675 66.075 ;
        RECT 138.125 64.885 138.295 65.055 ;
        RECT 139.965 65.225 140.135 65.395 ;
        RECT 140.425 65.565 140.595 65.735 ;
        RECT 141.805 65.905 141.975 66.075 ;
        RECT 140.885 64.885 141.055 65.055 ;
        RECT 144.565 65.905 144.735 66.075 ;
        RECT 145.945 65.905 146.115 66.075 ;
        RECT 145.025 65.565 145.195 65.735 ;
        RECT 143.645 64.885 143.815 65.055 ;
        RECT 145.945 64.885 146.115 65.055 ;
        RECT 91.205 64.375 91.375 64.545 ;
        RECT 91.665 64.375 91.835 64.545 ;
        RECT 92.125 64.375 92.295 64.545 ;
        RECT 92.585 64.375 92.755 64.545 ;
        RECT 93.045 64.375 93.215 64.545 ;
        RECT 93.505 64.375 93.675 64.545 ;
        RECT 93.965 64.375 94.135 64.545 ;
        RECT 94.425 64.375 94.595 64.545 ;
        RECT 94.885 64.375 95.055 64.545 ;
        RECT 95.345 64.375 95.515 64.545 ;
        RECT 95.805 64.375 95.975 64.545 ;
        RECT 96.265 64.375 96.435 64.545 ;
        RECT 96.725 64.375 96.895 64.545 ;
        RECT 97.185 64.375 97.355 64.545 ;
        RECT 97.645 64.375 97.815 64.545 ;
        RECT 98.105 64.375 98.275 64.545 ;
        RECT 98.565 64.375 98.735 64.545 ;
        RECT 99.025 64.375 99.195 64.545 ;
        RECT 99.485 64.375 99.655 64.545 ;
        RECT 99.945 64.375 100.115 64.545 ;
        RECT 100.405 64.375 100.575 64.545 ;
        RECT 100.865 64.375 101.035 64.545 ;
        RECT 101.325 64.375 101.495 64.545 ;
        RECT 101.785 64.375 101.955 64.545 ;
        RECT 102.245 64.375 102.415 64.545 ;
        RECT 102.705 64.375 102.875 64.545 ;
        RECT 103.165 64.375 103.335 64.545 ;
        RECT 103.625 64.375 103.795 64.545 ;
        RECT 104.085 64.375 104.255 64.545 ;
        RECT 104.545 64.375 104.715 64.545 ;
        RECT 105.005 64.375 105.175 64.545 ;
        RECT 105.465 64.375 105.635 64.545 ;
        RECT 105.925 64.375 106.095 64.545 ;
        RECT 106.385 64.375 106.555 64.545 ;
        RECT 106.845 64.375 107.015 64.545 ;
        RECT 107.305 64.375 107.475 64.545 ;
        RECT 107.765 64.375 107.935 64.545 ;
        RECT 108.225 64.375 108.395 64.545 ;
        RECT 108.685 64.375 108.855 64.545 ;
        RECT 109.145 64.375 109.315 64.545 ;
        RECT 109.605 64.375 109.775 64.545 ;
        RECT 110.065 64.375 110.235 64.545 ;
        RECT 110.525 64.375 110.695 64.545 ;
        RECT 110.985 64.375 111.155 64.545 ;
        RECT 111.445 64.375 111.615 64.545 ;
        RECT 111.905 64.375 112.075 64.545 ;
        RECT 112.365 64.375 112.535 64.545 ;
        RECT 112.825 64.375 112.995 64.545 ;
        RECT 113.285 64.375 113.455 64.545 ;
        RECT 113.745 64.375 113.915 64.545 ;
        RECT 114.205 64.375 114.375 64.545 ;
        RECT 114.665 64.375 114.835 64.545 ;
        RECT 115.125 64.375 115.295 64.545 ;
        RECT 115.585 64.375 115.755 64.545 ;
        RECT 116.045 64.375 116.215 64.545 ;
        RECT 116.505 64.375 116.675 64.545 ;
        RECT 116.965 64.375 117.135 64.545 ;
        RECT 117.425 64.375 117.595 64.545 ;
        RECT 117.885 64.375 118.055 64.545 ;
        RECT 118.345 64.375 118.515 64.545 ;
        RECT 118.805 64.375 118.975 64.545 ;
        RECT 119.265 64.375 119.435 64.545 ;
        RECT 119.725 64.375 119.895 64.545 ;
        RECT 120.185 64.375 120.355 64.545 ;
        RECT 120.645 64.375 120.815 64.545 ;
        RECT 121.105 64.375 121.275 64.545 ;
        RECT 121.565 64.375 121.735 64.545 ;
        RECT 122.025 64.375 122.195 64.545 ;
        RECT 122.485 64.375 122.655 64.545 ;
        RECT 122.945 64.375 123.115 64.545 ;
        RECT 123.405 64.375 123.575 64.545 ;
        RECT 123.865 64.375 124.035 64.545 ;
        RECT 124.325 64.375 124.495 64.545 ;
        RECT 124.785 64.375 124.955 64.545 ;
        RECT 125.245 64.375 125.415 64.545 ;
        RECT 125.705 64.375 125.875 64.545 ;
        RECT 126.165 64.375 126.335 64.545 ;
        RECT 126.625 64.375 126.795 64.545 ;
        RECT 127.085 64.375 127.255 64.545 ;
        RECT 127.545 64.375 127.715 64.545 ;
        RECT 128.005 64.375 128.175 64.545 ;
        RECT 128.465 64.375 128.635 64.545 ;
        RECT 128.925 64.375 129.095 64.545 ;
        RECT 129.385 64.375 129.555 64.545 ;
        RECT 129.845 64.375 130.015 64.545 ;
        RECT 130.305 64.375 130.475 64.545 ;
        RECT 130.765 64.375 130.935 64.545 ;
        RECT 131.225 64.375 131.395 64.545 ;
        RECT 131.685 64.375 131.855 64.545 ;
        RECT 132.145 64.375 132.315 64.545 ;
        RECT 132.605 64.375 132.775 64.545 ;
        RECT 133.065 64.375 133.235 64.545 ;
        RECT 133.525 64.375 133.695 64.545 ;
        RECT 133.985 64.375 134.155 64.545 ;
        RECT 134.445 64.375 134.615 64.545 ;
        RECT 134.905 64.375 135.075 64.545 ;
        RECT 135.365 64.375 135.535 64.545 ;
        RECT 135.825 64.375 135.995 64.545 ;
        RECT 136.285 64.375 136.455 64.545 ;
        RECT 136.745 64.375 136.915 64.545 ;
        RECT 137.205 64.375 137.375 64.545 ;
        RECT 137.665 64.375 137.835 64.545 ;
        RECT 138.125 64.375 138.295 64.545 ;
        RECT 138.585 64.375 138.755 64.545 ;
        RECT 139.045 64.375 139.215 64.545 ;
        RECT 139.505 64.375 139.675 64.545 ;
        RECT 139.965 64.375 140.135 64.545 ;
        RECT 140.425 64.375 140.595 64.545 ;
        RECT 140.885 64.375 141.055 64.545 ;
        RECT 141.345 64.375 141.515 64.545 ;
        RECT 141.805 64.375 141.975 64.545 ;
        RECT 142.265 64.375 142.435 64.545 ;
        RECT 142.725 64.375 142.895 64.545 ;
        RECT 143.185 64.375 143.355 64.545 ;
        RECT 143.645 64.375 143.815 64.545 ;
        RECT 144.105 64.375 144.275 64.545 ;
        RECT 144.565 64.375 144.735 64.545 ;
        RECT 145.025 64.375 145.195 64.545 ;
        RECT 145.485 64.375 145.655 64.545 ;
        RECT 145.945 64.375 146.115 64.545 ;
        RECT 146.405 64.375 146.575 64.545 ;
        RECT 146.865 64.375 147.035 64.545 ;
        RECT 147.325 64.375 147.495 64.545 ;
        RECT 147.785 64.375 147.955 64.545 ;
        RECT 148.245 64.375 148.415 64.545 ;
        RECT 148.705 64.375 148.875 64.545 ;
        RECT 149.165 64.375 149.335 64.545 ;
        RECT 149.625 64.375 149.795 64.545 ;
        RECT 150.085 64.375 150.255 64.545 ;
        RECT 150.545 64.375 150.715 64.545 ;
        RECT 151.005 64.375 151.175 64.545 ;
        RECT 151.465 64.375 151.635 64.545 ;
        RECT 151.925 64.375 152.095 64.545 ;
        RECT 95.905 63.525 96.075 63.695 ;
        RECT 93.045 62.165 93.215 62.335 ;
        RECT 94.825 62.820 94.995 62.990 ;
        RECT 94.525 62.505 94.695 62.675 ;
        RECT 95.905 62.845 96.075 63.015 ;
        RECT 99.025 63.525 99.195 63.695 ;
        RECT 97.765 62.505 97.935 62.675 ;
        RECT 98.125 62.505 98.295 62.675 ;
        RECT 99.485 62.845 99.655 63.015 ;
        RECT 100.915 63.525 101.085 63.695 ;
        RECT 100.405 62.505 100.575 62.675 ;
        RECT 101.320 62.845 101.490 63.015 ;
        RECT 101.785 63.185 101.955 63.355 ;
        RECT 103.165 62.845 103.335 63.015 ;
        RECT 102.705 62.165 102.875 62.335 ;
        RECT 106.720 63.185 106.890 63.355 ;
        RECT 105.925 62.165 106.095 62.335 ;
        RECT 107.765 62.845 107.935 63.015 ;
        RECT 107.305 62.165 107.475 62.335 ;
        RECT 109.145 62.845 109.315 63.015 ;
        RECT 110.525 63.525 110.695 63.695 ;
        RECT 109.605 62.165 109.775 62.335 ;
        RECT 112.825 62.845 112.995 63.015 ;
        RECT 113.290 62.845 113.460 63.015 ;
        RECT 111.905 62.505 112.075 62.675 ;
        RECT 113.695 63.525 113.865 63.695 ;
        RECT 114.205 62.505 114.375 62.675 ;
        RECT 115.585 63.525 115.755 63.695 ;
        RECT 115.125 62.845 115.295 63.015 ;
        RECT 118.705 63.525 118.875 63.695 ;
        RECT 116.845 62.505 117.015 62.675 ;
        RECT 118.705 62.845 118.875 63.015 ;
        RECT 119.785 62.820 119.955 62.990 ;
        RECT 120.085 62.505 120.255 62.675 ;
        RECT 121.565 62.165 121.735 62.335 ;
        RECT 122.025 62.165 122.195 62.335 ;
        RECT 127.085 63.865 127.255 64.035 ;
        RECT 124.785 62.845 124.955 63.015 ;
        RECT 126.625 62.845 126.795 63.015 ;
        RECT 142.265 62.845 142.435 63.015 ;
        RECT 143.185 62.845 143.355 63.015 ;
        RECT 142.725 62.165 142.895 62.335 ;
        RECT 146.865 63.865 147.035 64.035 ;
        RECT 147.325 62.845 147.495 63.015 ;
        RECT 32.720 61.595 32.890 61.765 ;
        RECT 91.205 61.655 91.375 61.825 ;
        RECT 91.665 61.655 91.835 61.825 ;
        RECT 92.125 61.655 92.295 61.825 ;
        RECT 92.585 61.655 92.755 61.825 ;
        RECT 93.045 61.655 93.215 61.825 ;
        RECT 93.505 61.655 93.675 61.825 ;
        RECT 93.965 61.655 94.135 61.825 ;
        RECT 94.425 61.655 94.595 61.825 ;
        RECT 94.885 61.655 95.055 61.825 ;
        RECT 95.345 61.655 95.515 61.825 ;
        RECT 95.805 61.655 95.975 61.825 ;
        RECT 96.265 61.655 96.435 61.825 ;
        RECT 96.725 61.655 96.895 61.825 ;
        RECT 97.185 61.655 97.355 61.825 ;
        RECT 97.645 61.655 97.815 61.825 ;
        RECT 98.105 61.655 98.275 61.825 ;
        RECT 98.565 61.655 98.735 61.825 ;
        RECT 99.025 61.655 99.195 61.825 ;
        RECT 99.485 61.655 99.655 61.825 ;
        RECT 99.945 61.655 100.115 61.825 ;
        RECT 100.405 61.655 100.575 61.825 ;
        RECT 100.865 61.655 101.035 61.825 ;
        RECT 101.325 61.655 101.495 61.825 ;
        RECT 101.785 61.655 101.955 61.825 ;
        RECT 102.245 61.655 102.415 61.825 ;
        RECT 102.705 61.655 102.875 61.825 ;
        RECT 103.165 61.655 103.335 61.825 ;
        RECT 103.625 61.655 103.795 61.825 ;
        RECT 104.085 61.655 104.255 61.825 ;
        RECT 104.545 61.655 104.715 61.825 ;
        RECT 105.005 61.655 105.175 61.825 ;
        RECT 105.465 61.655 105.635 61.825 ;
        RECT 105.925 61.655 106.095 61.825 ;
        RECT 106.385 61.655 106.555 61.825 ;
        RECT 106.845 61.655 107.015 61.825 ;
        RECT 107.305 61.655 107.475 61.825 ;
        RECT 107.765 61.655 107.935 61.825 ;
        RECT 108.225 61.655 108.395 61.825 ;
        RECT 108.685 61.655 108.855 61.825 ;
        RECT 109.145 61.655 109.315 61.825 ;
        RECT 109.605 61.655 109.775 61.825 ;
        RECT 110.065 61.655 110.235 61.825 ;
        RECT 110.525 61.655 110.695 61.825 ;
        RECT 110.985 61.655 111.155 61.825 ;
        RECT 111.445 61.655 111.615 61.825 ;
        RECT 111.905 61.655 112.075 61.825 ;
        RECT 112.365 61.655 112.535 61.825 ;
        RECT 112.825 61.655 112.995 61.825 ;
        RECT 113.285 61.655 113.455 61.825 ;
        RECT 113.745 61.655 113.915 61.825 ;
        RECT 114.205 61.655 114.375 61.825 ;
        RECT 114.665 61.655 114.835 61.825 ;
        RECT 115.125 61.655 115.295 61.825 ;
        RECT 115.585 61.655 115.755 61.825 ;
        RECT 116.045 61.655 116.215 61.825 ;
        RECT 116.505 61.655 116.675 61.825 ;
        RECT 116.965 61.655 117.135 61.825 ;
        RECT 117.425 61.655 117.595 61.825 ;
        RECT 117.885 61.655 118.055 61.825 ;
        RECT 118.345 61.655 118.515 61.825 ;
        RECT 118.805 61.655 118.975 61.825 ;
        RECT 119.265 61.655 119.435 61.825 ;
        RECT 119.725 61.655 119.895 61.825 ;
        RECT 120.185 61.655 120.355 61.825 ;
        RECT 120.645 61.655 120.815 61.825 ;
        RECT 121.105 61.655 121.275 61.825 ;
        RECT 121.565 61.655 121.735 61.825 ;
        RECT 122.025 61.655 122.195 61.825 ;
        RECT 122.485 61.655 122.655 61.825 ;
        RECT 122.945 61.655 123.115 61.825 ;
        RECT 123.405 61.655 123.575 61.825 ;
        RECT 123.865 61.655 124.035 61.825 ;
        RECT 124.325 61.655 124.495 61.825 ;
        RECT 124.785 61.655 124.955 61.825 ;
        RECT 125.245 61.655 125.415 61.825 ;
        RECT 125.705 61.655 125.875 61.825 ;
        RECT 126.165 61.655 126.335 61.825 ;
        RECT 126.625 61.655 126.795 61.825 ;
        RECT 127.085 61.655 127.255 61.825 ;
        RECT 127.545 61.655 127.715 61.825 ;
        RECT 128.005 61.655 128.175 61.825 ;
        RECT 128.465 61.655 128.635 61.825 ;
        RECT 128.925 61.655 129.095 61.825 ;
        RECT 129.385 61.655 129.555 61.825 ;
        RECT 129.845 61.655 130.015 61.825 ;
        RECT 130.305 61.655 130.475 61.825 ;
        RECT 130.765 61.655 130.935 61.825 ;
        RECT 131.225 61.655 131.395 61.825 ;
        RECT 131.685 61.655 131.855 61.825 ;
        RECT 132.145 61.655 132.315 61.825 ;
        RECT 132.605 61.655 132.775 61.825 ;
        RECT 133.065 61.655 133.235 61.825 ;
        RECT 133.525 61.655 133.695 61.825 ;
        RECT 133.985 61.655 134.155 61.825 ;
        RECT 134.445 61.655 134.615 61.825 ;
        RECT 134.905 61.655 135.075 61.825 ;
        RECT 135.365 61.655 135.535 61.825 ;
        RECT 135.825 61.655 135.995 61.825 ;
        RECT 136.285 61.655 136.455 61.825 ;
        RECT 136.745 61.655 136.915 61.825 ;
        RECT 137.205 61.655 137.375 61.825 ;
        RECT 137.665 61.655 137.835 61.825 ;
        RECT 138.125 61.655 138.295 61.825 ;
        RECT 138.585 61.655 138.755 61.825 ;
        RECT 139.045 61.655 139.215 61.825 ;
        RECT 139.505 61.655 139.675 61.825 ;
        RECT 139.965 61.655 140.135 61.825 ;
        RECT 140.425 61.655 140.595 61.825 ;
        RECT 140.885 61.655 141.055 61.825 ;
        RECT 141.345 61.655 141.515 61.825 ;
        RECT 141.805 61.655 141.975 61.825 ;
        RECT 142.265 61.655 142.435 61.825 ;
        RECT 142.725 61.655 142.895 61.825 ;
        RECT 143.185 61.655 143.355 61.825 ;
        RECT 143.645 61.655 143.815 61.825 ;
        RECT 144.105 61.655 144.275 61.825 ;
        RECT 144.565 61.655 144.735 61.825 ;
        RECT 145.025 61.655 145.195 61.825 ;
        RECT 145.485 61.655 145.655 61.825 ;
        RECT 145.945 61.655 146.115 61.825 ;
        RECT 146.405 61.655 146.575 61.825 ;
        RECT 146.865 61.655 147.035 61.825 ;
        RECT 147.325 61.655 147.495 61.825 ;
        RECT 147.785 61.655 147.955 61.825 ;
        RECT 148.245 61.655 148.415 61.825 ;
        RECT 148.705 61.655 148.875 61.825 ;
        RECT 149.165 61.655 149.335 61.825 ;
        RECT 149.625 61.655 149.795 61.825 ;
        RECT 150.085 61.655 150.255 61.825 ;
        RECT 150.545 61.655 150.715 61.825 ;
        RECT 151.005 61.655 151.175 61.825 ;
        RECT 151.465 61.655 151.635 61.825 ;
        RECT 151.925 61.655 152.095 61.825 ;
        RECT 97.645 60.805 97.815 60.975 ;
        RECT 97.185 60.465 97.355 60.635 ;
        RECT 98.105 60.465 98.275 60.635 ;
        RECT 98.565 60.465 98.735 60.635 ;
        RECT 29.875 59.300 30.055 59.475 ;
        RECT 101.785 61.145 101.955 61.315 ;
        RECT 99.485 60.465 99.655 60.635 ;
        RECT 99.945 60.465 100.115 60.635 ;
        RECT 100.405 60.465 100.575 60.635 ;
        RECT 102.245 61.145 102.415 61.315 ;
        RECT 103.165 60.805 103.335 60.975 ;
        RECT 105.465 60.805 105.635 60.975 ;
        RECT 103.165 59.445 103.335 59.615 ;
        RECT 105.005 59.785 105.175 59.955 ;
        RECT 114.205 61.145 114.375 61.315 ;
        RECT 106.385 60.465 106.555 60.635 ;
        RECT 107.305 60.465 107.475 60.635 ;
        RECT 107.765 60.465 107.935 60.635 ;
        RECT 116.045 61.145 116.215 61.315 ;
        RECT 117.425 60.805 117.595 60.975 ;
        RECT 115.125 60.465 115.295 60.635 ;
        RECT 116.505 60.465 116.675 60.635 ;
        RECT 123.865 59.445 124.035 59.615 ;
        RECT 145.945 60.465 146.115 60.635 ;
        RECT 147.325 60.805 147.495 60.975 ;
        RECT 146.405 59.785 146.575 59.955 ;
        RECT 91.205 58.935 91.375 59.105 ;
        RECT 91.665 58.935 91.835 59.105 ;
        RECT 92.125 58.935 92.295 59.105 ;
        RECT 92.585 58.935 92.755 59.105 ;
        RECT 93.045 58.935 93.215 59.105 ;
        RECT 93.505 58.935 93.675 59.105 ;
        RECT 93.965 58.935 94.135 59.105 ;
        RECT 94.425 58.935 94.595 59.105 ;
        RECT 94.885 58.935 95.055 59.105 ;
        RECT 95.345 58.935 95.515 59.105 ;
        RECT 95.805 58.935 95.975 59.105 ;
        RECT 96.265 58.935 96.435 59.105 ;
        RECT 96.725 58.935 96.895 59.105 ;
        RECT 97.185 58.935 97.355 59.105 ;
        RECT 97.645 58.935 97.815 59.105 ;
        RECT 98.105 58.935 98.275 59.105 ;
        RECT 98.565 58.935 98.735 59.105 ;
        RECT 99.025 58.935 99.195 59.105 ;
        RECT 99.485 58.935 99.655 59.105 ;
        RECT 99.945 58.935 100.115 59.105 ;
        RECT 100.405 58.935 100.575 59.105 ;
        RECT 100.865 58.935 101.035 59.105 ;
        RECT 101.325 58.935 101.495 59.105 ;
        RECT 101.785 58.935 101.955 59.105 ;
        RECT 102.245 58.935 102.415 59.105 ;
        RECT 102.705 58.935 102.875 59.105 ;
        RECT 103.165 58.935 103.335 59.105 ;
        RECT 103.625 58.935 103.795 59.105 ;
        RECT 104.085 58.935 104.255 59.105 ;
        RECT 104.545 58.935 104.715 59.105 ;
        RECT 105.005 58.935 105.175 59.105 ;
        RECT 105.465 58.935 105.635 59.105 ;
        RECT 105.925 58.935 106.095 59.105 ;
        RECT 106.385 58.935 106.555 59.105 ;
        RECT 106.845 58.935 107.015 59.105 ;
        RECT 107.305 58.935 107.475 59.105 ;
        RECT 107.765 58.935 107.935 59.105 ;
        RECT 108.225 58.935 108.395 59.105 ;
        RECT 108.685 58.935 108.855 59.105 ;
        RECT 109.145 58.935 109.315 59.105 ;
        RECT 109.605 58.935 109.775 59.105 ;
        RECT 110.065 58.935 110.235 59.105 ;
        RECT 110.525 58.935 110.695 59.105 ;
        RECT 110.985 58.935 111.155 59.105 ;
        RECT 111.445 58.935 111.615 59.105 ;
        RECT 111.905 58.935 112.075 59.105 ;
        RECT 112.365 58.935 112.535 59.105 ;
        RECT 112.825 58.935 112.995 59.105 ;
        RECT 113.285 58.935 113.455 59.105 ;
        RECT 113.745 58.935 113.915 59.105 ;
        RECT 114.205 58.935 114.375 59.105 ;
        RECT 114.665 58.935 114.835 59.105 ;
        RECT 115.125 58.935 115.295 59.105 ;
        RECT 115.585 58.935 115.755 59.105 ;
        RECT 116.045 58.935 116.215 59.105 ;
        RECT 116.505 58.935 116.675 59.105 ;
        RECT 116.965 58.935 117.135 59.105 ;
        RECT 117.425 58.935 117.595 59.105 ;
        RECT 117.885 58.935 118.055 59.105 ;
        RECT 118.345 58.935 118.515 59.105 ;
        RECT 118.805 58.935 118.975 59.105 ;
        RECT 119.265 58.935 119.435 59.105 ;
        RECT 119.725 58.935 119.895 59.105 ;
        RECT 120.185 58.935 120.355 59.105 ;
        RECT 120.645 58.935 120.815 59.105 ;
        RECT 121.105 58.935 121.275 59.105 ;
        RECT 121.565 58.935 121.735 59.105 ;
        RECT 122.025 58.935 122.195 59.105 ;
        RECT 122.485 58.935 122.655 59.105 ;
        RECT 122.945 58.935 123.115 59.105 ;
        RECT 123.405 58.935 123.575 59.105 ;
        RECT 123.865 58.935 124.035 59.105 ;
        RECT 124.325 58.935 124.495 59.105 ;
        RECT 124.785 58.935 124.955 59.105 ;
        RECT 125.245 58.935 125.415 59.105 ;
        RECT 125.705 58.935 125.875 59.105 ;
        RECT 126.165 58.935 126.335 59.105 ;
        RECT 126.625 58.935 126.795 59.105 ;
        RECT 127.085 58.935 127.255 59.105 ;
        RECT 127.545 58.935 127.715 59.105 ;
        RECT 128.005 58.935 128.175 59.105 ;
        RECT 128.465 58.935 128.635 59.105 ;
        RECT 128.925 58.935 129.095 59.105 ;
        RECT 129.385 58.935 129.555 59.105 ;
        RECT 129.845 58.935 130.015 59.105 ;
        RECT 130.305 58.935 130.475 59.105 ;
        RECT 130.765 58.935 130.935 59.105 ;
        RECT 131.225 58.935 131.395 59.105 ;
        RECT 131.685 58.935 131.855 59.105 ;
        RECT 132.145 58.935 132.315 59.105 ;
        RECT 132.605 58.935 132.775 59.105 ;
        RECT 133.065 58.935 133.235 59.105 ;
        RECT 133.525 58.935 133.695 59.105 ;
        RECT 133.985 58.935 134.155 59.105 ;
        RECT 134.445 58.935 134.615 59.105 ;
        RECT 134.905 58.935 135.075 59.105 ;
        RECT 135.365 58.935 135.535 59.105 ;
        RECT 135.825 58.935 135.995 59.105 ;
        RECT 136.285 58.935 136.455 59.105 ;
        RECT 136.745 58.935 136.915 59.105 ;
        RECT 137.205 58.935 137.375 59.105 ;
        RECT 137.665 58.935 137.835 59.105 ;
        RECT 138.125 58.935 138.295 59.105 ;
        RECT 138.585 58.935 138.755 59.105 ;
        RECT 139.045 58.935 139.215 59.105 ;
        RECT 139.505 58.935 139.675 59.105 ;
        RECT 139.965 58.935 140.135 59.105 ;
        RECT 140.425 58.935 140.595 59.105 ;
        RECT 140.885 58.935 141.055 59.105 ;
        RECT 141.345 58.935 141.515 59.105 ;
        RECT 141.805 58.935 141.975 59.105 ;
        RECT 142.265 58.935 142.435 59.105 ;
        RECT 142.725 58.935 142.895 59.105 ;
        RECT 143.185 58.935 143.355 59.105 ;
        RECT 143.645 58.935 143.815 59.105 ;
        RECT 144.105 58.935 144.275 59.105 ;
        RECT 144.565 58.935 144.735 59.105 ;
        RECT 145.025 58.935 145.195 59.105 ;
        RECT 145.485 58.935 145.655 59.105 ;
        RECT 145.945 58.935 146.115 59.105 ;
        RECT 146.405 58.935 146.575 59.105 ;
        RECT 146.865 58.935 147.035 59.105 ;
        RECT 147.325 58.935 147.495 59.105 ;
        RECT 147.785 58.935 147.955 59.105 ;
        RECT 148.245 58.935 148.415 59.105 ;
        RECT 148.705 58.935 148.875 59.105 ;
        RECT 149.165 58.935 149.335 59.105 ;
        RECT 149.625 58.935 149.795 59.105 ;
        RECT 150.085 58.935 150.255 59.105 ;
        RECT 150.545 58.935 150.715 59.105 ;
        RECT 151.005 58.935 151.175 59.105 ;
        RECT 151.465 58.935 151.635 59.105 ;
        RECT 151.925 58.935 152.095 59.105 ;
        RECT 26.535 57.930 26.900 58.460 ;
        RECT 23.180 56.600 23.630 57.180 ;
        RECT 96.725 57.745 96.895 57.915 ;
        RECT 98.565 58.425 98.735 58.595 ;
        RECT 97.645 57.405 97.815 57.575 ;
        RECT 98.105 57.405 98.275 57.575 ;
        RECT 100.865 58.425 101.035 58.595 ;
        RECT 99.485 57.405 99.655 57.575 ;
        RECT 100.405 57.405 100.575 57.575 ;
        RECT 101.785 57.405 101.955 57.575 ;
        RECT 102.245 57.405 102.415 57.575 ;
        RECT 113.285 58.425 113.455 58.595 ;
        RECT 120.645 57.405 120.815 57.575 ;
        RECT 126.165 57.405 126.335 57.575 ;
        RECT 126.625 57.405 126.795 57.575 ;
        RECT 125.705 56.725 125.875 56.895 ;
        RECT 127.545 56.725 127.715 56.895 ;
        RECT 132.145 57.745 132.315 57.915 ;
        RECT 131.225 57.065 131.395 57.235 ;
        RECT 133.985 57.405 134.155 57.575 ;
        RECT 133.065 56.725 133.235 56.895 ;
        RECT 141.345 57.405 141.515 57.575 ;
        RECT 141.810 57.405 141.980 57.575 ;
        RECT 142.215 58.085 142.385 58.255 ;
        RECT 142.725 57.745 142.895 57.915 ;
        RECT 144.105 58.085 144.275 58.255 ;
        RECT 143.645 57.405 143.815 57.575 ;
        RECT 147.225 58.085 147.395 58.255 ;
        RECT 145.365 57.065 145.535 57.235 ;
        RECT 147.225 57.405 147.395 57.575 ;
        RECT 150.085 58.425 150.255 58.595 ;
        RECT 148.305 57.380 148.475 57.550 ;
        RECT 148.605 57.065 148.775 57.235 ;
        RECT 91.205 56.215 91.375 56.385 ;
        RECT 91.665 56.215 91.835 56.385 ;
        RECT 92.125 56.215 92.295 56.385 ;
        RECT 92.585 56.215 92.755 56.385 ;
        RECT 93.045 56.215 93.215 56.385 ;
        RECT 93.505 56.215 93.675 56.385 ;
        RECT 93.965 56.215 94.135 56.385 ;
        RECT 94.425 56.215 94.595 56.385 ;
        RECT 94.885 56.215 95.055 56.385 ;
        RECT 95.345 56.215 95.515 56.385 ;
        RECT 95.805 56.215 95.975 56.385 ;
        RECT 96.265 56.215 96.435 56.385 ;
        RECT 96.725 56.215 96.895 56.385 ;
        RECT 97.185 56.215 97.355 56.385 ;
        RECT 97.645 56.215 97.815 56.385 ;
        RECT 98.105 56.215 98.275 56.385 ;
        RECT 98.565 56.215 98.735 56.385 ;
        RECT 99.025 56.215 99.195 56.385 ;
        RECT 99.485 56.215 99.655 56.385 ;
        RECT 99.945 56.215 100.115 56.385 ;
        RECT 100.405 56.215 100.575 56.385 ;
        RECT 100.865 56.215 101.035 56.385 ;
        RECT 101.325 56.215 101.495 56.385 ;
        RECT 101.785 56.215 101.955 56.385 ;
        RECT 102.245 56.215 102.415 56.385 ;
        RECT 102.705 56.215 102.875 56.385 ;
        RECT 103.165 56.215 103.335 56.385 ;
        RECT 103.625 56.215 103.795 56.385 ;
        RECT 104.085 56.215 104.255 56.385 ;
        RECT 104.545 56.215 104.715 56.385 ;
        RECT 105.005 56.215 105.175 56.385 ;
        RECT 105.465 56.215 105.635 56.385 ;
        RECT 105.925 56.215 106.095 56.385 ;
        RECT 106.385 56.215 106.555 56.385 ;
        RECT 106.845 56.215 107.015 56.385 ;
        RECT 107.305 56.215 107.475 56.385 ;
        RECT 107.765 56.215 107.935 56.385 ;
        RECT 108.225 56.215 108.395 56.385 ;
        RECT 108.685 56.215 108.855 56.385 ;
        RECT 109.145 56.215 109.315 56.385 ;
        RECT 109.605 56.215 109.775 56.385 ;
        RECT 110.065 56.215 110.235 56.385 ;
        RECT 110.525 56.215 110.695 56.385 ;
        RECT 110.985 56.215 111.155 56.385 ;
        RECT 111.445 56.215 111.615 56.385 ;
        RECT 111.905 56.215 112.075 56.385 ;
        RECT 112.365 56.215 112.535 56.385 ;
        RECT 112.825 56.215 112.995 56.385 ;
        RECT 113.285 56.215 113.455 56.385 ;
        RECT 113.745 56.215 113.915 56.385 ;
        RECT 114.205 56.215 114.375 56.385 ;
        RECT 114.665 56.215 114.835 56.385 ;
        RECT 115.125 56.215 115.295 56.385 ;
        RECT 115.585 56.215 115.755 56.385 ;
        RECT 116.045 56.215 116.215 56.385 ;
        RECT 116.505 56.215 116.675 56.385 ;
        RECT 116.965 56.215 117.135 56.385 ;
        RECT 117.425 56.215 117.595 56.385 ;
        RECT 117.885 56.215 118.055 56.385 ;
        RECT 118.345 56.215 118.515 56.385 ;
        RECT 118.805 56.215 118.975 56.385 ;
        RECT 119.265 56.215 119.435 56.385 ;
        RECT 119.725 56.215 119.895 56.385 ;
        RECT 120.185 56.215 120.355 56.385 ;
        RECT 120.645 56.215 120.815 56.385 ;
        RECT 121.105 56.215 121.275 56.385 ;
        RECT 121.565 56.215 121.735 56.385 ;
        RECT 122.025 56.215 122.195 56.385 ;
        RECT 122.485 56.215 122.655 56.385 ;
        RECT 122.945 56.215 123.115 56.385 ;
        RECT 123.405 56.215 123.575 56.385 ;
        RECT 123.865 56.215 124.035 56.385 ;
        RECT 124.325 56.215 124.495 56.385 ;
        RECT 124.785 56.215 124.955 56.385 ;
        RECT 125.245 56.215 125.415 56.385 ;
        RECT 125.705 56.215 125.875 56.385 ;
        RECT 126.165 56.215 126.335 56.385 ;
        RECT 126.625 56.215 126.795 56.385 ;
        RECT 127.085 56.215 127.255 56.385 ;
        RECT 127.545 56.215 127.715 56.385 ;
        RECT 128.005 56.215 128.175 56.385 ;
        RECT 128.465 56.215 128.635 56.385 ;
        RECT 128.925 56.215 129.095 56.385 ;
        RECT 129.385 56.215 129.555 56.385 ;
        RECT 129.845 56.215 130.015 56.385 ;
        RECT 130.305 56.215 130.475 56.385 ;
        RECT 130.765 56.215 130.935 56.385 ;
        RECT 131.225 56.215 131.395 56.385 ;
        RECT 131.685 56.215 131.855 56.385 ;
        RECT 132.145 56.215 132.315 56.385 ;
        RECT 132.605 56.215 132.775 56.385 ;
        RECT 133.065 56.215 133.235 56.385 ;
        RECT 133.525 56.215 133.695 56.385 ;
        RECT 133.985 56.215 134.155 56.385 ;
        RECT 134.445 56.215 134.615 56.385 ;
        RECT 134.905 56.215 135.075 56.385 ;
        RECT 135.365 56.215 135.535 56.385 ;
        RECT 135.825 56.215 135.995 56.385 ;
        RECT 136.285 56.215 136.455 56.385 ;
        RECT 136.745 56.215 136.915 56.385 ;
        RECT 137.205 56.215 137.375 56.385 ;
        RECT 137.665 56.215 137.835 56.385 ;
        RECT 138.125 56.215 138.295 56.385 ;
        RECT 138.585 56.215 138.755 56.385 ;
        RECT 139.045 56.215 139.215 56.385 ;
        RECT 139.505 56.215 139.675 56.385 ;
        RECT 139.965 56.215 140.135 56.385 ;
        RECT 140.425 56.215 140.595 56.385 ;
        RECT 140.885 56.215 141.055 56.385 ;
        RECT 141.345 56.215 141.515 56.385 ;
        RECT 141.805 56.215 141.975 56.385 ;
        RECT 142.265 56.215 142.435 56.385 ;
        RECT 142.725 56.215 142.895 56.385 ;
        RECT 143.185 56.215 143.355 56.385 ;
        RECT 143.645 56.215 143.815 56.385 ;
        RECT 144.105 56.215 144.275 56.385 ;
        RECT 144.565 56.215 144.735 56.385 ;
        RECT 145.025 56.215 145.195 56.385 ;
        RECT 145.485 56.215 145.655 56.385 ;
        RECT 145.945 56.215 146.115 56.385 ;
        RECT 146.405 56.215 146.575 56.385 ;
        RECT 146.865 56.215 147.035 56.385 ;
        RECT 147.325 56.215 147.495 56.385 ;
        RECT 147.785 56.215 147.955 56.385 ;
        RECT 148.245 56.215 148.415 56.385 ;
        RECT 148.705 56.215 148.875 56.385 ;
        RECT 149.165 56.215 149.335 56.385 ;
        RECT 149.625 56.215 149.795 56.385 ;
        RECT 150.085 56.215 150.255 56.385 ;
        RECT 150.545 56.215 150.715 56.385 ;
        RECT 151.005 56.215 151.175 56.385 ;
        RECT 151.465 56.215 151.635 56.385 ;
        RECT 151.925 56.215 152.095 56.385 ;
        RECT 6.110 53.600 6.300 55.585 ;
        RECT 99.025 55.705 99.195 55.875 ;
        RECT 98.565 55.025 98.735 55.195 ;
        RECT 99.485 55.025 99.655 55.195 ;
        RECT 112.365 54.345 112.535 54.515 ;
        RECT 115.125 55.705 115.295 55.875 ;
        RECT 114.205 55.365 114.375 55.535 ;
        RECT 114.205 54.005 114.375 54.175 ;
        RECT 116.505 55.025 116.675 55.195 ;
        RECT 118.345 55.025 118.515 55.195 ;
        RECT 115.585 54.005 115.755 54.175 ;
        RECT 118.805 54.005 118.975 54.175 ;
        RECT 123.505 55.365 123.675 55.535 ;
        RECT 123.805 55.050 123.975 55.220 ;
        RECT 122.025 54.005 122.195 54.175 ;
        RECT 124.885 55.025 125.055 55.195 ;
        RECT 126.745 55.365 126.915 55.535 ;
        RECT 127.105 55.365 127.275 55.535 ;
        RECT 124.885 54.345 125.055 54.515 ;
        RECT 128.465 55.025 128.635 55.195 ;
        RECT 128.005 54.345 128.175 54.515 ;
        RECT 129.385 55.365 129.555 55.535 ;
        RECT 129.895 54.345 130.065 54.515 ;
        RECT 130.300 55.025 130.470 55.195 ;
        RECT 130.765 55.025 130.935 55.195 ;
        RECT 131.685 55.025 131.855 55.195 ;
        RECT 132.150 55.025 132.320 55.195 ;
        RECT 133.065 55.365 133.235 55.535 ;
        RECT 132.555 54.345 132.725 54.515 ;
        RECT 133.985 55.025 134.155 55.195 ;
        RECT 135.345 55.365 135.515 55.535 ;
        RECT 135.705 55.365 135.875 55.535 ;
        RECT 134.445 54.345 134.615 54.515 ;
        RECT 137.565 55.025 137.735 55.195 ;
        RECT 138.945 55.365 139.115 55.535 ;
        RECT 138.645 55.050 138.815 55.220 ;
        RECT 137.565 54.345 137.735 54.515 ;
        RECT 141.805 55.025 141.975 55.195 ;
        RECT 140.425 54.005 140.595 54.175 ;
        RECT 141.345 54.685 141.515 54.855 ;
        RECT 146.405 55.025 146.575 55.195 ;
        RECT 146.865 54.005 147.035 54.175 ;
        RECT 91.205 53.495 91.375 53.665 ;
        RECT 91.665 53.495 91.835 53.665 ;
        RECT 92.125 53.495 92.295 53.665 ;
        RECT 92.585 53.495 92.755 53.665 ;
        RECT 93.045 53.495 93.215 53.665 ;
        RECT 93.505 53.495 93.675 53.665 ;
        RECT 93.965 53.495 94.135 53.665 ;
        RECT 94.425 53.495 94.595 53.665 ;
        RECT 94.885 53.495 95.055 53.665 ;
        RECT 95.345 53.495 95.515 53.665 ;
        RECT 95.805 53.495 95.975 53.665 ;
        RECT 96.265 53.495 96.435 53.665 ;
        RECT 96.725 53.495 96.895 53.665 ;
        RECT 97.185 53.495 97.355 53.665 ;
        RECT 97.645 53.495 97.815 53.665 ;
        RECT 98.105 53.495 98.275 53.665 ;
        RECT 98.565 53.495 98.735 53.665 ;
        RECT 99.025 53.495 99.195 53.665 ;
        RECT 99.485 53.495 99.655 53.665 ;
        RECT 99.945 53.495 100.115 53.665 ;
        RECT 100.405 53.495 100.575 53.665 ;
        RECT 100.865 53.495 101.035 53.665 ;
        RECT 101.325 53.495 101.495 53.665 ;
        RECT 101.785 53.495 101.955 53.665 ;
        RECT 102.245 53.495 102.415 53.665 ;
        RECT 102.705 53.495 102.875 53.665 ;
        RECT 103.165 53.495 103.335 53.665 ;
        RECT 103.625 53.495 103.795 53.665 ;
        RECT 104.085 53.495 104.255 53.665 ;
        RECT 104.545 53.495 104.715 53.665 ;
        RECT 105.005 53.495 105.175 53.665 ;
        RECT 105.465 53.495 105.635 53.665 ;
        RECT 105.925 53.495 106.095 53.665 ;
        RECT 106.385 53.495 106.555 53.665 ;
        RECT 106.845 53.495 107.015 53.665 ;
        RECT 107.305 53.495 107.475 53.665 ;
        RECT 107.765 53.495 107.935 53.665 ;
        RECT 108.225 53.495 108.395 53.665 ;
        RECT 108.685 53.495 108.855 53.665 ;
        RECT 109.145 53.495 109.315 53.665 ;
        RECT 109.605 53.495 109.775 53.665 ;
        RECT 110.065 53.495 110.235 53.665 ;
        RECT 110.525 53.495 110.695 53.665 ;
        RECT 110.985 53.495 111.155 53.665 ;
        RECT 111.445 53.495 111.615 53.665 ;
        RECT 111.905 53.495 112.075 53.665 ;
        RECT 112.365 53.495 112.535 53.665 ;
        RECT 112.825 53.495 112.995 53.665 ;
        RECT 113.285 53.495 113.455 53.665 ;
        RECT 113.745 53.495 113.915 53.665 ;
        RECT 114.205 53.495 114.375 53.665 ;
        RECT 114.665 53.495 114.835 53.665 ;
        RECT 115.125 53.495 115.295 53.665 ;
        RECT 115.585 53.495 115.755 53.665 ;
        RECT 116.045 53.495 116.215 53.665 ;
        RECT 116.505 53.495 116.675 53.665 ;
        RECT 116.965 53.495 117.135 53.665 ;
        RECT 117.425 53.495 117.595 53.665 ;
        RECT 117.885 53.495 118.055 53.665 ;
        RECT 118.345 53.495 118.515 53.665 ;
        RECT 118.805 53.495 118.975 53.665 ;
        RECT 119.265 53.495 119.435 53.665 ;
        RECT 119.725 53.495 119.895 53.665 ;
        RECT 120.185 53.495 120.355 53.665 ;
        RECT 120.645 53.495 120.815 53.665 ;
        RECT 121.105 53.495 121.275 53.665 ;
        RECT 121.565 53.495 121.735 53.665 ;
        RECT 122.025 53.495 122.195 53.665 ;
        RECT 122.485 53.495 122.655 53.665 ;
        RECT 122.945 53.495 123.115 53.665 ;
        RECT 123.405 53.495 123.575 53.665 ;
        RECT 123.865 53.495 124.035 53.665 ;
        RECT 124.325 53.495 124.495 53.665 ;
        RECT 124.785 53.495 124.955 53.665 ;
        RECT 125.245 53.495 125.415 53.665 ;
        RECT 125.705 53.495 125.875 53.665 ;
        RECT 126.165 53.495 126.335 53.665 ;
        RECT 126.625 53.495 126.795 53.665 ;
        RECT 127.085 53.495 127.255 53.665 ;
        RECT 127.545 53.495 127.715 53.665 ;
        RECT 128.005 53.495 128.175 53.665 ;
        RECT 128.465 53.495 128.635 53.665 ;
        RECT 128.925 53.495 129.095 53.665 ;
        RECT 129.385 53.495 129.555 53.665 ;
        RECT 129.845 53.495 130.015 53.665 ;
        RECT 130.305 53.495 130.475 53.665 ;
        RECT 130.765 53.495 130.935 53.665 ;
        RECT 131.225 53.495 131.395 53.665 ;
        RECT 131.685 53.495 131.855 53.665 ;
        RECT 132.145 53.495 132.315 53.665 ;
        RECT 132.605 53.495 132.775 53.665 ;
        RECT 133.065 53.495 133.235 53.665 ;
        RECT 133.525 53.495 133.695 53.665 ;
        RECT 133.985 53.495 134.155 53.665 ;
        RECT 134.445 53.495 134.615 53.665 ;
        RECT 134.905 53.495 135.075 53.665 ;
        RECT 135.365 53.495 135.535 53.665 ;
        RECT 135.825 53.495 135.995 53.665 ;
        RECT 136.285 53.495 136.455 53.665 ;
        RECT 136.745 53.495 136.915 53.665 ;
        RECT 137.205 53.495 137.375 53.665 ;
        RECT 137.665 53.495 137.835 53.665 ;
        RECT 138.125 53.495 138.295 53.665 ;
        RECT 138.585 53.495 138.755 53.665 ;
        RECT 139.045 53.495 139.215 53.665 ;
        RECT 139.505 53.495 139.675 53.665 ;
        RECT 139.965 53.495 140.135 53.665 ;
        RECT 140.425 53.495 140.595 53.665 ;
        RECT 140.885 53.495 141.055 53.665 ;
        RECT 141.345 53.495 141.515 53.665 ;
        RECT 141.805 53.495 141.975 53.665 ;
        RECT 142.265 53.495 142.435 53.665 ;
        RECT 142.725 53.495 142.895 53.665 ;
        RECT 143.185 53.495 143.355 53.665 ;
        RECT 143.645 53.495 143.815 53.665 ;
        RECT 144.105 53.495 144.275 53.665 ;
        RECT 144.565 53.495 144.735 53.665 ;
        RECT 145.025 53.495 145.195 53.665 ;
        RECT 145.485 53.495 145.655 53.665 ;
        RECT 145.945 53.495 146.115 53.665 ;
        RECT 146.405 53.495 146.575 53.665 ;
        RECT 146.865 53.495 147.035 53.665 ;
        RECT 147.325 53.495 147.495 53.665 ;
        RECT 147.785 53.495 147.955 53.665 ;
        RECT 148.245 53.495 148.415 53.665 ;
        RECT 148.705 53.495 148.875 53.665 ;
        RECT 149.165 53.495 149.335 53.665 ;
        RECT 149.625 53.495 149.795 53.665 ;
        RECT 150.085 53.495 150.255 53.665 ;
        RECT 150.545 53.495 150.715 53.665 ;
        RECT 151.005 53.495 151.175 53.665 ;
        RECT 151.465 53.495 151.635 53.665 ;
        RECT 151.925 53.495 152.095 53.665 ;
        RECT 6.100 51.015 6.300 51.245 ;
        RECT 92.585 51.965 92.755 52.135 ;
        RECT 93.050 51.965 93.220 52.135 ;
        RECT 93.455 52.645 93.625 52.815 ;
        RECT 93.900 52.985 94.070 53.155 ;
        RECT 95.345 52.645 95.515 52.815 ;
        RECT 94.885 51.965 95.055 52.135 ;
        RECT 98.465 52.645 98.635 52.815 ;
        RECT 96.605 51.625 96.775 51.795 ;
        RECT 98.465 51.965 98.635 52.135 ;
        RECT 99.545 51.940 99.715 52.110 ;
        RECT 99.845 51.625 100.015 51.795 ;
        RECT 102.705 51.965 102.875 52.135 ;
        RECT 101.325 51.285 101.495 51.455 ;
        RECT 102.245 51.625 102.415 51.795 ;
        RECT 107.305 51.625 107.475 51.795 ;
        RECT 108.225 51.285 108.395 51.455 ;
        RECT 110.065 51.965 110.235 52.135 ;
        RECT 109.145 51.285 109.315 51.455 ;
        RECT 111.905 51.625 112.075 51.795 ;
        RECT 113.285 52.305 113.455 52.475 ;
        RECT 113.750 51.965 113.920 52.135 ;
        RECT 112.825 51.625 112.995 51.795 ;
        RECT 114.155 52.645 114.325 52.815 ;
        RECT 114.600 52.985 114.770 53.155 ;
        RECT 116.045 52.645 116.215 52.815 ;
        RECT 115.585 51.965 115.755 52.135 ;
        RECT 119.165 52.645 119.335 52.815 ;
        RECT 117.305 51.625 117.475 51.795 ;
        RECT 119.165 51.965 119.335 52.135 ;
        RECT 120.245 51.940 120.415 52.110 ;
        RECT 120.545 51.625 120.715 51.795 ;
        RECT 123.405 51.965 123.575 52.135 ;
        RECT 124.325 51.965 124.495 52.135 ;
        RECT 125.245 51.965 125.415 52.135 ;
        RECT 122.025 51.285 122.195 51.455 ;
        RECT 125.705 51.965 125.875 52.135 ;
        RECT 127.545 52.985 127.715 53.155 ;
        RECT 128.465 52.985 128.635 53.155 ;
        RECT 132.145 52.985 132.315 53.155 ;
        RECT 131.225 52.645 131.395 52.815 ;
        RECT 127.545 51.285 127.715 51.455 ;
        RECT 132.145 51.625 132.315 51.795 ;
        RECT 133.985 51.965 134.155 52.135 ;
        RECT 135.365 52.985 135.535 53.155 ;
        RECT 134.445 51.285 134.615 51.455 ;
        RECT 135.285 51.285 135.455 51.455 ;
        RECT 136.745 51.965 136.915 52.135 ;
        RECT 138.585 52.985 138.755 53.155 ;
        RECT 136.285 51.625 136.455 51.795 ;
        RECT 139.965 51.965 140.135 52.135 ;
        RECT 138.585 51.285 138.755 51.455 ;
        RECT 139.505 51.285 139.675 51.455 ;
        RECT 141.345 51.965 141.515 52.135 ;
        RECT 141.810 51.965 141.980 52.135 ;
        RECT 140.885 51.285 141.055 51.455 ;
        RECT 142.215 52.645 142.385 52.815 ;
        RECT 142.725 51.625 142.895 51.795 ;
        RECT 144.105 52.645 144.275 52.815 ;
        RECT 143.645 51.965 143.815 52.135 ;
        RECT 147.225 52.645 147.395 52.815 ;
        RECT 145.365 51.625 145.535 51.795 ;
        RECT 147.225 51.965 147.395 52.135 ;
        RECT 150.085 52.305 150.255 52.475 ;
        RECT 148.305 51.940 148.475 52.110 ;
        RECT 148.605 51.625 148.775 51.795 ;
        RECT 91.205 50.775 91.375 50.945 ;
        RECT 91.665 50.775 91.835 50.945 ;
        RECT 92.125 50.775 92.295 50.945 ;
        RECT 92.585 50.775 92.755 50.945 ;
        RECT 93.045 50.775 93.215 50.945 ;
        RECT 93.505 50.775 93.675 50.945 ;
        RECT 93.965 50.775 94.135 50.945 ;
        RECT 94.425 50.775 94.595 50.945 ;
        RECT 94.885 50.775 95.055 50.945 ;
        RECT 95.345 50.775 95.515 50.945 ;
        RECT 95.805 50.775 95.975 50.945 ;
        RECT 96.265 50.775 96.435 50.945 ;
        RECT 96.725 50.775 96.895 50.945 ;
        RECT 97.185 50.775 97.355 50.945 ;
        RECT 97.645 50.775 97.815 50.945 ;
        RECT 98.105 50.775 98.275 50.945 ;
        RECT 98.565 50.775 98.735 50.945 ;
        RECT 99.025 50.775 99.195 50.945 ;
        RECT 99.485 50.775 99.655 50.945 ;
        RECT 99.945 50.775 100.115 50.945 ;
        RECT 100.405 50.775 100.575 50.945 ;
        RECT 100.865 50.775 101.035 50.945 ;
        RECT 101.325 50.775 101.495 50.945 ;
        RECT 101.785 50.775 101.955 50.945 ;
        RECT 102.245 50.775 102.415 50.945 ;
        RECT 102.705 50.775 102.875 50.945 ;
        RECT 103.165 50.775 103.335 50.945 ;
        RECT 103.625 50.775 103.795 50.945 ;
        RECT 104.085 50.775 104.255 50.945 ;
        RECT 104.545 50.775 104.715 50.945 ;
        RECT 105.005 50.775 105.175 50.945 ;
        RECT 105.465 50.775 105.635 50.945 ;
        RECT 105.925 50.775 106.095 50.945 ;
        RECT 106.385 50.775 106.555 50.945 ;
        RECT 106.845 50.775 107.015 50.945 ;
        RECT 107.305 50.775 107.475 50.945 ;
        RECT 107.765 50.775 107.935 50.945 ;
        RECT 108.225 50.775 108.395 50.945 ;
        RECT 108.685 50.775 108.855 50.945 ;
        RECT 109.145 50.775 109.315 50.945 ;
        RECT 109.605 50.775 109.775 50.945 ;
        RECT 110.065 50.775 110.235 50.945 ;
        RECT 110.525 50.775 110.695 50.945 ;
        RECT 110.985 50.775 111.155 50.945 ;
        RECT 111.445 50.775 111.615 50.945 ;
        RECT 111.905 50.775 112.075 50.945 ;
        RECT 112.365 50.775 112.535 50.945 ;
        RECT 112.825 50.775 112.995 50.945 ;
        RECT 113.285 50.775 113.455 50.945 ;
        RECT 113.745 50.775 113.915 50.945 ;
        RECT 114.205 50.775 114.375 50.945 ;
        RECT 114.665 50.775 114.835 50.945 ;
        RECT 115.125 50.775 115.295 50.945 ;
        RECT 115.585 50.775 115.755 50.945 ;
        RECT 116.045 50.775 116.215 50.945 ;
        RECT 116.505 50.775 116.675 50.945 ;
        RECT 116.965 50.775 117.135 50.945 ;
        RECT 117.425 50.775 117.595 50.945 ;
        RECT 117.885 50.775 118.055 50.945 ;
        RECT 118.345 50.775 118.515 50.945 ;
        RECT 118.805 50.775 118.975 50.945 ;
        RECT 119.265 50.775 119.435 50.945 ;
        RECT 119.725 50.775 119.895 50.945 ;
        RECT 120.185 50.775 120.355 50.945 ;
        RECT 120.645 50.775 120.815 50.945 ;
        RECT 121.105 50.775 121.275 50.945 ;
        RECT 121.565 50.775 121.735 50.945 ;
        RECT 122.025 50.775 122.195 50.945 ;
        RECT 122.485 50.775 122.655 50.945 ;
        RECT 122.945 50.775 123.115 50.945 ;
        RECT 123.405 50.775 123.575 50.945 ;
        RECT 123.865 50.775 124.035 50.945 ;
        RECT 124.325 50.775 124.495 50.945 ;
        RECT 124.785 50.775 124.955 50.945 ;
        RECT 125.245 50.775 125.415 50.945 ;
        RECT 125.705 50.775 125.875 50.945 ;
        RECT 126.165 50.775 126.335 50.945 ;
        RECT 126.625 50.775 126.795 50.945 ;
        RECT 127.085 50.775 127.255 50.945 ;
        RECT 127.545 50.775 127.715 50.945 ;
        RECT 128.005 50.775 128.175 50.945 ;
        RECT 128.465 50.775 128.635 50.945 ;
        RECT 128.925 50.775 129.095 50.945 ;
        RECT 129.385 50.775 129.555 50.945 ;
        RECT 129.845 50.775 130.015 50.945 ;
        RECT 130.305 50.775 130.475 50.945 ;
        RECT 130.765 50.775 130.935 50.945 ;
        RECT 131.225 50.775 131.395 50.945 ;
        RECT 131.685 50.775 131.855 50.945 ;
        RECT 132.145 50.775 132.315 50.945 ;
        RECT 132.605 50.775 132.775 50.945 ;
        RECT 133.065 50.775 133.235 50.945 ;
        RECT 133.525 50.775 133.695 50.945 ;
        RECT 133.985 50.775 134.155 50.945 ;
        RECT 134.445 50.775 134.615 50.945 ;
        RECT 134.905 50.775 135.075 50.945 ;
        RECT 135.365 50.775 135.535 50.945 ;
        RECT 135.825 50.775 135.995 50.945 ;
        RECT 136.285 50.775 136.455 50.945 ;
        RECT 136.745 50.775 136.915 50.945 ;
        RECT 137.205 50.775 137.375 50.945 ;
        RECT 137.665 50.775 137.835 50.945 ;
        RECT 138.125 50.775 138.295 50.945 ;
        RECT 138.585 50.775 138.755 50.945 ;
        RECT 139.045 50.775 139.215 50.945 ;
        RECT 139.505 50.775 139.675 50.945 ;
        RECT 139.965 50.775 140.135 50.945 ;
        RECT 140.425 50.775 140.595 50.945 ;
        RECT 140.885 50.775 141.055 50.945 ;
        RECT 141.345 50.775 141.515 50.945 ;
        RECT 141.805 50.775 141.975 50.945 ;
        RECT 142.265 50.775 142.435 50.945 ;
        RECT 142.725 50.775 142.895 50.945 ;
        RECT 143.185 50.775 143.355 50.945 ;
        RECT 143.645 50.775 143.815 50.945 ;
        RECT 144.105 50.775 144.275 50.945 ;
        RECT 144.565 50.775 144.735 50.945 ;
        RECT 145.025 50.775 145.195 50.945 ;
        RECT 145.485 50.775 145.655 50.945 ;
        RECT 145.945 50.775 146.115 50.945 ;
        RECT 146.405 50.775 146.575 50.945 ;
        RECT 146.865 50.775 147.035 50.945 ;
        RECT 147.325 50.775 147.495 50.945 ;
        RECT 147.785 50.775 147.955 50.945 ;
        RECT 148.245 50.775 148.415 50.945 ;
        RECT 148.705 50.775 148.875 50.945 ;
        RECT 149.165 50.775 149.335 50.945 ;
        RECT 149.625 50.775 149.795 50.945 ;
        RECT 150.085 50.775 150.255 50.945 ;
        RECT 150.545 50.775 150.715 50.945 ;
        RECT 151.005 50.775 151.175 50.945 ;
        RECT 151.465 50.775 151.635 50.945 ;
        RECT 151.925 50.775 152.095 50.945 ;
        RECT 98.565 49.585 98.735 49.755 ;
        RECT 99.945 49.585 100.115 49.755 ;
        RECT 97.645 48.565 97.815 48.735 ;
        RECT 99.485 48.565 99.655 48.735 ;
        RECT 103.165 49.585 103.335 49.755 ;
        RECT 102.245 49.245 102.415 49.415 ;
        RECT 104.085 49.245 104.255 49.415 ;
        RECT 105.005 50.265 105.175 50.435 ;
        RECT 105.695 49.755 105.865 49.925 ;
        RECT 106.845 49.925 107.015 50.095 ;
        RECT 107.305 49.585 107.475 49.755 ;
        RECT 107.770 49.585 107.940 49.755 ;
        RECT 108.685 49.925 108.855 50.095 ;
        RECT 108.175 48.905 108.345 49.075 ;
        RECT 105.925 48.565 106.095 48.735 ;
        RECT 109.605 49.585 109.775 49.755 ;
        RECT 110.965 49.925 111.135 50.095 ;
        RECT 111.325 49.925 111.495 50.095 ;
        RECT 110.065 48.905 110.235 49.075 ;
        RECT 113.185 49.585 113.355 49.755 ;
        RECT 114.565 49.925 114.735 50.095 ;
        RECT 114.265 49.610 114.435 49.780 ;
        RECT 113.185 48.905 113.355 49.075 ;
        RECT 116.045 49.245 116.215 49.415 ;
        RECT 128.465 50.265 128.635 50.435 ;
        RECT 126.625 49.585 126.795 49.755 ;
        RECT 127.545 49.585 127.715 49.755 ;
        RECT 132.145 49.245 132.315 49.415 ;
        RECT 133.065 49.925 133.235 50.095 ;
        RECT 133.525 49.585 133.695 49.755 ;
        RECT 133.985 50.265 134.155 50.435 ;
        RECT 137.205 50.265 137.375 50.435 ;
        RECT 134.905 49.925 135.075 50.095 ;
        RECT 135.365 49.925 135.535 50.095 ;
        RECT 136.285 49.925 136.455 50.095 ;
        RECT 149.165 49.585 149.335 49.755 ;
        RECT 150.545 49.245 150.715 49.415 ;
        RECT 91.205 48.055 91.375 48.225 ;
        RECT 91.665 48.055 91.835 48.225 ;
        RECT 92.125 48.055 92.295 48.225 ;
        RECT 92.585 48.055 92.755 48.225 ;
        RECT 93.045 48.055 93.215 48.225 ;
        RECT 93.505 48.055 93.675 48.225 ;
        RECT 93.965 48.055 94.135 48.225 ;
        RECT 94.425 48.055 94.595 48.225 ;
        RECT 94.885 48.055 95.055 48.225 ;
        RECT 95.345 48.055 95.515 48.225 ;
        RECT 95.805 48.055 95.975 48.225 ;
        RECT 96.265 48.055 96.435 48.225 ;
        RECT 96.725 48.055 96.895 48.225 ;
        RECT 97.185 48.055 97.355 48.225 ;
        RECT 97.645 48.055 97.815 48.225 ;
        RECT 98.105 48.055 98.275 48.225 ;
        RECT 98.565 48.055 98.735 48.225 ;
        RECT 99.025 48.055 99.195 48.225 ;
        RECT 99.485 48.055 99.655 48.225 ;
        RECT 99.945 48.055 100.115 48.225 ;
        RECT 100.405 48.055 100.575 48.225 ;
        RECT 100.865 48.055 101.035 48.225 ;
        RECT 101.325 48.055 101.495 48.225 ;
        RECT 101.785 48.055 101.955 48.225 ;
        RECT 102.245 48.055 102.415 48.225 ;
        RECT 102.705 48.055 102.875 48.225 ;
        RECT 103.165 48.055 103.335 48.225 ;
        RECT 103.625 48.055 103.795 48.225 ;
        RECT 104.085 48.055 104.255 48.225 ;
        RECT 104.545 48.055 104.715 48.225 ;
        RECT 105.005 48.055 105.175 48.225 ;
        RECT 105.465 48.055 105.635 48.225 ;
        RECT 105.925 48.055 106.095 48.225 ;
        RECT 106.385 48.055 106.555 48.225 ;
        RECT 106.845 48.055 107.015 48.225 ;
        RECT 107.305 48.055 107.475 48.225 ;
        RECT 107.765 48.055 107.935 48.225 ;
        RECT 108.225 48.055 108.395 48.225 ;
        RECT 108.685 48.055 108.855 48.225 ;
        RECT 109.145 48.055 109.315 48.225 ;
        RECT 109.605 48.055 109.775 48.225 ;
        RECT 110.065 48.055 110.235 48.225 ;
        RECT 110.525 48.055 110.695 48.225 ;
        RECT 110.985 48.055 111.155 48.225 ;
        RECT 111.445 48.055 111.615 48.225 ;
        RECT 111.905 48.055 112.075 48.225 ;
        RECT 112.365 48.055 112.535 48.225 ;
        RECT 112.825 48.055 112.995 48.225 ;
        RECT 113.285 48.055 113.455 48.225 ;
        RECT 113.745 48.055 113.915 48.225 ;
        RECT 114.205 48.055 114.375 48.225 ;
        RECT 114.665 48.055 114.835 48.225 ;
        RECT 115.125 48.055 115.295 48.225 ;
        RECT 115.585 48.055 115.755 48.225 ;
        RECT 116.045 48.055 116.215 48.225 ;
        RECT 116.505 48.055 116.675 48.225 ;
        RECT 116.965 48.055 117.135 48.225 ;
        RECT 117.425 48.055 117.595 48.225 ;
        RECT 117.885 48.055 118.055 48.225 ;
        RECT 118.345 48.055 118.515 48.225 ;
        RECT 118.805 48.055 118.975 48.225 ;
        RECT 119.265 48.055 119.435 48.225 ;
        RECT 119.725 48.055 119.895 48.225 ;
        RECT 120.185 48.055 120.355 48.225 ;
        RECT 120.645 48.055 120.815 48.225 ;
        RECT 121.105 48.055 121.275 48.225 ;
        RECT 121.565 48.055 121.735 48.225 ;
        RECT 122.025 48.055 122.195 48.225 ;
        RECT 122.485 48.055 122.655 48.225 ;
        RECT 122.945 48.055 123.115 48.225 ;
        RECT 123.405 48.055 123.575 48.225 ;
        RECT 123.865 48.055 124.035 48.225 ;
        RECT 124.325 48.055 124.495 48.225 ;
        RECT 124.785 48.055 124.955 48.225 ;
        RECT 125.245 48.055 125.415 48.225 ;
        RECT 125.705 48.055 125.875 48.225 ;
        RECT 126.165 48.055 126.335 48.225 ;
        RECT 126.625 48.055 126.795 48.225 ;
        RECT 127.085 48.055 127.255 48.225 ;
        RECT 127.545 48.055 127.715 48.225 ;
        RECT 128.005 48.055 128.175 48.225 ;
        RECT 128.465 48.055 128.635 48.225 ;
        RECT 128.925 48.055 129.095 48.225 ;
        RECT 129.385 48.055 129.555 48.225 ;
        RECT 129.845 48.055 130.015 48.225 ;
        RECT 130.305 48.055 130.475 48.225 ;
        RECT 130.765 48.055 130.935 48.225 ;
        RECT 131.225 48.055 131.395 48.225 ;
        RECT 131.685 48.055 131.855 48.225 ;
        RECT 132.145 48.055 132.315 48.225 ;
        RECT 132.605 48.055 132.775 48.225 ;
        RECT 133.065 48.055 133.235 48.225 ;
        RECT 133.525 48.055 133.695 48.225 ;
        RECT 133.985 48.055 134.155 48.225 ;
        RECT 134.445 48.055 134.615 48.225 ;
        RECT 134.905 48.055 135.075 48.225 ;
        RECT 135.365 48.055 135.535 48.225 ;
        RECT 135.825 48.055 135.995 48.225 ;
        RECT 136.285 48.055 136.455 48.225 ;
        RECT 136.745 48.055 136.915 48.225 ;
        RECT 137.205 48.055 137.375 48.225 ;
        RECT 137.665 48.055 137.835 48.225 ;
        RECT 138.125 48.055 138.295 48.225 ;
        RECT 138.585 48.055 138.755 48.225 ;
        RECT 139.045 48.055 139.215 48.225 ;
        RECT 139.505 48.055 139.675 48.225 ;
        RECT 139.965 48.055 140.135 48.225 ;
        RECT 140.425 48.055 140.595 48.225 ;
        RECT 140.885 48.055 141.055 48.225 ;
        RECT 141.345 48.055 141.515 48.225 ;
        RECT 141.805 48.055 141.975 48.225 ;
        RECT 142.265 48.055 142.435 48.225 ;
        RECT 142.725 48.055 142.895 48.225 ;
        RECT 143.185 48.055 143.355 48.225 ;
        RECT 143.645 48.055 143.815 48.225 ;
        RECT 144.105 48.055 144.275 48.225 ;
        RECT 144.565 48.055 144.735 48.225 ;
        RECT 145.025 48.055 145.195 48.225 ;
        RECT 145.485 48.055 145.655 48.225 ;
        RECT 145.945 48.055 146.115 48.225 ;
        RECT 146.405 48.055 146.575 48.225 ;
        RECT 146.865 48.055 147.035 48.225 ;
        RECT 147.325 48.055 147.495 48.225 ;
        RECT 147.785 48.055 147.955 48.225 ;
        RECT 148.245 48.055 148.415 48.225 ;
        RECT 148.705 48.055 148.875 48.225 ;
        RECT 149.165 48.055 149.335 48.225 ;
        RECT 149.625 48.055 149.795 48.225 ;
        RECT 150.085 48.055 150.255 48.225 ;
        RECT 150.545 48.055 150.715 48.225 ;
        RECT 151.005 48.055 151.175 48.225 ;
        RECT 151.465 48.055 151.635 48.225 ;
        RECT 151.925 48.055 152.095 48.225 ;
        RECT 6.110 44.505 6.300 46.490 ;
        RECT 93.045 46.865 93.215 47.035 ;
        RECT 93.510 46.525 93.680 46.695 ;
        RECT 93.915 47.205 94.085 47.375 ;
        RECT 94.425 46.865 94.595 47.035 ;
        RECT 95.805 47.205 95.975 47.375 ;
        RECT 95.345 46.525 95.515 46.695 ;
        RECT 98.925 47.205 99.095 47.375 ;
        RECT 97.065 46.185 97.235 46.355 ;
        RECT 98.925 46.525 99.095 46.695 ;
        RECT 100.005 46.500 100.175 46.670 ;
        RECT 100.305 46.185 100.475 46.355 ;
        RECT 101.785 45.845 101.955 46.015 ;
        RECT 105.465 47.205 105.635 47.375 ;
        RECT 107.305 47.545 107.475 47.715 ;
        RECT 107.305 46.185 107.475 46.355 ;
        RECT 110.985 47.545 111.155 47.715 ;
        RECT 117.885 47.545 118.055 47.715 ;
        RECT 108.225 45.845 108.395 46.015 ;
        RECT 117.425 46.185 117.595 46.355 ;
        RECT 120.745 47.205 120.915 47.375 ;
        RECT 119.665 46.500 119.835 46.670 ;
        RECT 119.365 46.185 119.535 46.355 ;
        RECT 120.745 46.525 120.915 46.695 ;
        RECT 123.865 47.205 124.035 47.375 ;
        RECT 122.605 46.185 122.775 46.355 ;
        RECT 122.965 46.185 123.135 46.355 ;
        RECT 124.325 46.525 124.495 46.695 ;
        RECT 125.755 47.205 125.925 47.375 ;
        RECT 125.245 46.865 125.415 47.035 ;
        RECT 126.160 46.525 126.330 46.695 ;
        RECT 126.625 46.865 126.795 47.035 ;
        RECT 127.085 46.525 127.255 46.695 ;
        RECT 127.545 46.185 127.715 46.355 ;
        RECT 91.205 45.335 91.375 45.505 ;
        RECT 91.665 45.335 91.835 45.505 ;
        RECT 92.125 45.335 92.295 45.505 ;
        RECT 92.585 45.335 92.755 45.505 ;
        RECT 93.045 45.335 93.215 45.505 ;
        RECT 93.505 45.335 93.675 45.505 ;
        RECT 93.965 45.335 94.135 45.505 ;
        RECT 94.425 45.335 94.595 45.505 ;
        RECT 94.885 45.335 95.055 45.505 ;
        RECT 95.345 45.335 95.515 45.505 ;
        RECT 95.805 45.335 95.975 45.505 ;
        RECT 96.265 45.335 96.435 45.505 ;
        RECT 96.725 45.335 96.895 45.505 ;
        RECT 97.185 45.335 97.355 45.505 ;
        RECT 97.645 45.335 97.815 45.505 ;
        RECT 98.105 45.335 98.275 45.505 ;
        RECT 98.565 45.335 98.735 45.505 ;
        RECT 99.025 45.335 99.195 45.505 ;
        RECT 99.485 45.335 99.655 45.505 ;
        RECT 99.945 45.335 100.115 45.505 ;
        RECT 100.405 45.335 100.575 45.505 ;
        RECT 100.865 45.335 101.035 45.505 ;
        RECT 101.325 45.335 101.495 45.505 ;
        RECT 101.785 45.335 101.955 45.505 ;
        RECT 102.245 45.335 102.415 45.505 ;
        RECT 102.705 45.335 102.875 45.505 ;
        RECT 103.165 45.335 103.335 45.505 ;
        RECT 103.625 45.335 103.795 45.505 ;
        RECT 104.085 45.335 104.255 45.505 ;
        RECT 104.545 45.335 104.715 45.505 ;
        RECT 105.005 45.335 105.175 45.505 ;
        RECT 105.465 45.335 105.635 45.505 ;
        RECT 105.925 45.335 106.095 45.505 ;
        RECT 106.385 45.335 106.555 45.505 ;
        RECT 106.845 45.335 107.015 45.505 ;
        RECT 107.305 45.335 107.475 45.505 ;
        RECT 107.765 45.335 107.935 45.505 ;
        RECT 108.225 45.335 108.395 45.505 ;
        RECT 108.685 45.335 108.855 45.505 ;
        RECT 109.145 45.335 109.315 45.505 ;
        RECT 109.605 45.335 109.775 45.505 ;
        RECT 110.065 45.335 110.235 45.505 ;
        RECT 110.525 45.335 110.695 45.505 ;
        RECT 110.985 45.335 111.155 45.505 ;
        RECT 111.445 45.335 111.615 45.505 ;
        RECT 111.905 45.335 112.075 45.505 ;
        RECT 112.365 45.335 112.535 45.505 ;
        RECT 112.825 45.335 112.995 45.505 ;
        RECT 113.285 45.335 113.455 45.505 ;
        RECT 113.745 45.335 113.915 45.505 ;
        RECT 114.205 45.335 114.375 45.505 ;
        RECT 114.665 45.335 114.835 45.505 ;
        RECT 115.125 45.335 115.295 45.505 ;
        RECT 115.585 45.335 115.755 45.505 ;
        RECT 116.045 45.335 116.215 45.505 ;
        RECT 116.505 45.335 116.675 45.505 ;
        RECT 116.965 45.335 117.135 45.505 ;
        RECT 117.425 45.335 117.595 45.505 ;
        RECT 117.885 45.335 118.055 45.505 ;
        RECT 118.345 45.335 118.515 45.505 ;
        RECT 118.805 45.335 118.975 45.505 ;
        RECT 119.265 45.335 119.435 45.505 ;
        RECT 119.725 45.335 119.895 45.505 ;
        RECT 120.185 45.335 120.355 45.505 ;
        RECT 120.645 45.335 120.815 45.505 ;
        RECT 121.105 45.335 121.275 45.505 ;
        RECT 121.565 45.335 121.735 45.505 ;
        RECT 122.025 45.335 122.195 45.505 ;
        RECT 122.485 45.335 122.655 45.505 ;
        RECT 122.945 45.335 123.115 45.505 ;
        RECT 123.405 45.335 123.575 45.505 ;
        RECT 123.865 45.335 124.035 45.505 ;
        RECT 124.325 45.335 124.495 45.505 ;
        RECT 124.785 45.335 124.955 45.505 ;
        RECT 125.245 45.335 125.415 45.505 ;
        RECT 125.705 45.335 125.875 45.505 ;
        RECT 126.165 45.335 126.335 45.505 ;
        RECT 126.625 45.335 126.795 45.505 ;
        RECT 127.085 45.335 127.255 45.505 ;
        RECT 127.545 45.335 127.715 45.505 ;
        RECT 128.005 45.335 128.175 45.505 ;
        RECT 128.465 45.335 128.635 45.505 ;
        RECT 128.925 45.335 129.095 45.505 ;
        RECT 129.385 45.335 129.555 45.505 ;
        RECT 129.845 45.335 130.015 45.505 ;
        RECT 130.305 45.335 130.475 45.505 ;
        RECT 130.765 45.335 130.935 45.505 ;
        RECT 131.225 45.335 131.395 45.505 ;
        RECT 131.685 45.335 131.855 45.505 ;
        RECT 132.145 45.335 132.315 45.505 ;
        RECT 132.605 45.335 132.775 45.505 ;
        RECT 133.065 45.335 133.235 45.505 ;
        RECT 133.525 45.335 133.695 45.505 ;
        RECT 133.985 45.335 134.155 45.505 ;
        RECT 134.445 45.335 134.615 45.505 ;
        RECT 134.905 45.335 135.075 45.505 ;
        RECT 135.365 45.335 135.535 45.505 ;
        RECT 135.825 45.335 135.995 45.505 ;
        RECT 136.285 45.335 136.455 45.505 ;
        RECT 136.745 45.335 136.915 45.505 ;
        RECT 137.205 45.335 137.375 45.505 ;
        RECT 137.665 45.335 137.835 45.505 ;
        RECT 138.125 45.335 138.295 45.505 ;
        RECT 138.585 45.335 138.755 45.505 ;
        RECT 139.045 45.335 139.215 45.505 ;
        RECT 139.505 45.335 139.675 45.505 ;
        RECT 139.965 45.335 140.135 45.505 ;
        RECT 140.425 45.335 140.595 45.505 ;
        RECT 140.885 45.335 141.055 45.505 ;
        RECT 141.345 45.335 141.515 45.505 ;
        RECT 141.805 45.335 141.975 45.505 ;
        RECT 142.265 45.335 142.435 45.505 ;
        RECT 142.725 45.335 142.895 45.505 ;
        RECT 143.185 45.335 143.355 45.505 ;
        RECT 143.645 45.335 143.815 45.505 ;
        RECT 144.105 45.335 144.275 45.505 ;
        RECT 144.565 45.335 144.735 45.505 ;
        RECT 145.025 45.335 145.195 45.505 ;
        RECT 145.485 45.335 145.655 45.505 ;
        RECT 145.945 45.335 146.115 45.505 ;
        RECT 146.405 45.335 146.575 45.505 ;
        RECT 146.865 45.335 147.035 45.505 ;
        RECT 147.325 45.335 147.495 45.505 ;
        RECT 147.785 45.335 147.955 45.505 ;
        RECT 148.245 45.335 148.415 45.505 ;
        RECT 148.705 45.335 148.875 45.505 ;
        RECT 149.165 45.335 149.335 45.505 ;
        RECT 149.625 45.335 149.795 45.505 ;
        RECT 150.085 45.335 150.255 45.505 ;
        RECT 150.545 45.335 150.715 45.505 ;
        RECT 151.005 45.335 151.175 45.505 ;
        RECT 151.465 45.335 151.635 45.505 ;
        RECT 151.925 45.335 152.095 45.505 ;
        RECT 99.485 44.825 99.655 44.995 ;
        RECT 96.265 44.145 96.435 44.315 ;
        RECT 6.110 41.350 6.300 43.335 ;
        RECT 100.405 44.485 100.575 44.655 ;
        RECT 100.405 43.125 100.575 43.295 ;
        RECT 102.245 44.145 102.415 44.315 ;
        RECT 104.545 44.485 104.715 44.655 ;
        RECT 105.465 44.145 105.635 44.315 ;
        RECT 106.385 44.485 106.555 44.655 ;
        RECT 110.525 44.825 110.695 44.995 ;
        RECT 111.445 44.485 111.615 44.655 ;
        RECT 111.905 44.145 112.075 44.315 ;
        RECT 112.365 44.825 112.535 44.995 ;
        RECT 113.285 44.485 113.455 44.655 ;
        RECT 114.205 44.825 114.375 44.995 ;
        RECT 114.665 44.145 114.835 44.315 ;
        RECT 122.485 44.145 122.655 44.315 ;
        RECT 129.385 44.825 129.555 44.995 ;
        RECT 126.955 44.485 127.125 44.655 ;
        RECT 127.545 44.145 127.715 44.315 ;
        RECT 128.005 44.145 128.175 44.315 ;
        RECT 128.465 44.145 128.635 44.315 ;
        RECT 125.705 43.805 125.875 43.975 ;
        RECT 132.145 44.145 132.315 44.315 ;
        RECT 134.445 44.145 134.615 44.315 ;
        RECT 137.665 44.825 137.835 44.995 ;
        RECT 131.685 43.125 131.855 43.295 ;
        RECT 133.985 43.125 134.155 43.295 ;
        RECT 136.745 44.145 136.915 44.315 ;
        RECT 138.125 44.485 138.295 44.655 ;
        RECT 137.665 44.145 137.835 44.315 ;
        RECT 139.045 44.485 139.215 44.655 ;
        RECT 140.425 44.485 140.595 44.655 ;
        RECT 142.265 44.825 142.435 44.995 ;
        RECT 141.425 44.485 141.595 44.655 ;
        RECT 139.965 43.125 140.135 43.295 ;
        RECT 141.345 43.125 141.515 43.295 ;
        RECT 144.105 44.145 144.275 44.315 ;
        RECT 146.405 44.145 146.575 44.315 ;
        RECT 143.185 43.125 143.355 43.295 ;
        RECT 146.865 43.125 147.035 43.295 ;
        RECT 91.205 42.615 91.375 42.785 ;
        RECT 91.665 42.615 91.835 42.785 ;
        RECT 92.125 42.615 92.295 42.785 ;
        RECT 92.585 42.615 92.755 42.785 ;
        RECT 93.045 42.615 93.215 42.785 ;
        RECT 93.505 42.615 93.675 42.785 ;
        RECT 93.965 42.615 94.135 42.785 ;
        RECT 94.425 42.615 94.595 42.785 ;
        RECT 94.885 42.615 95.055 42.785 ;
        RECT 95.345 42.615 95.515 42.785 ;
        RECT 95.805 42.615 95.975 42.785 ;
        RECT 96.265 42.615 96.435 42.785 ;
        RECT 96.725 42.615 96.895 42.785 ;
        RECT 97.185 42.615 97.355 42.785 ;
        RECT 97.645 42.615 97.815 42.785 ;
        RECT 98.105 42.615 98.275 42.785 ;
        RECT 98.565 42.615 98.735 42.785 ;
        RECT 99.025 42.615 99.195 42.785 ;
        RECT 99.485 42.615 99.655 42.785 ;
        RECT 99.945 42.615 100.115 42.785 ;
        RECT 100.405 42.615 100.575 42.785 ;
        RECT 100.865 42.615 101.035 42.785 ;
        RECT 101.325 42.615 101.495 42.785 ;
        RECT 101.785 42.615 101.955 42.785 ;
        RECT 102.245 42.615 102.415 42.785 ;
        RECT 102.705 42.615 102.875 42.785 ;
        RECT 103.165 42.615 103.335 42.785 ;
        RECT 103.625 42.615 103.795 42.785 ;
        RECT 104.085 42.615 104.255 42.785 ;
        RECT 104.545 42.615 104.715 42.785 ;
        RECT 105.005 42.615 105.175 42.785 ;
        RECT 105.465 42.615 105.635 42.785 ;
        RECT 105.925 42.615 106.095 42.785 ;
        RECT 106.385 42.615 106.555 42.785 ;
        RECT 106.845 42.615 107.015 42.785 ;
        RECT 107.305 42.615 107.475 42.785 ;
        RECT 107.765 42.615 107.935 42.785 ;
        RECT 108.225 42.615 108.395 42.785 ;
        RECT 108.685 42.615 108.855 42.785 ;
        RECT 109.145 42.615 109.315 42.785 ;
        RECT 109.605 42.615 109.775 42.785 ;
        RECT 110.065 42.615 110.235 42.785 ;
        RECT 110.525 42.615 110.695 42.785 ;
        RECT 110.985 42.615 111.155 42.785 ;
        RECT 111.445 42.615 111.615 42.785 ;
        RECT 111.905 42.615 112.075 42.785 ;
        RECT 112.365 42.615 112.535 42.785 ;
        RECT 112.825 42.615 112.995 42.785 ;
        RECT 113.285 42.615 113.455 42.785 ;
        RECT 113.745 42.615 113.915 42.785 ;
        RECT 114.205 42.615 114.375 42.785 ;
        RECT 114.665 42.615 114.835 42.785 ;
        RECT 115.125 42.615 115.295 42.785 ;
        RECT 115.585 42.615 115.755 42.785 ;
        RECT 116.045 42.615 116.215 42.785 ;
        RECT 116.505 42.615 116.675 42.785 ;
        RECT 116.965 42.615 117.135 42.785 ;
        RECT 117.425 42.615 117.595 42.785 ;
        RECT 117.885 42.615 118.055 42.785 ;
        RECT 118.345 42.615 118.515 42.785 ;
        RECT 118.805 42.615 118.975 42.785 ;
        RECT 119.265 42.615 119.435 42.785 ;
        RECT 119.725 42.615 119.895 42.785 ;
        RECT 120.185 42.615 120.355 42.785 ;
        RECT 120.645 42.615 120.815 42.785 ;
        RECT 121.105 42.615 121.275 42.785 ;
        RECT 121.565 42.615 121.735 42.785 ;
        RECT 122.025 42.615 122.195 42.785 ;
        RECT 122.485 42.615 122.655 42.785 ;
        RECT 122.945 42.615 123.115 42.785 ;
        RECT 123.405 42.615 123.575 42.785 ;
        RECT 123.865 42.615 124.035 42.785 ;
        RECT 124.325 42.615 124.495 42.785 ;
        RECT 124.785 42.615 124.955 42.785 ;
        RECT 125.245 42.615 125.415 42.785 ;
        RECT 125.705 42.615 125.875 42.785 ;
        RECT 126.165 42.615 126.335 42.785 ;
        RECT 126.625 42.615 126.795 42.785 ;
        RECT 127.085 42.615 127.255 42.785 ;
        RECT 127.545 42.615 127.715 42.785 ;
        RECT 128.005 42.615 128.175 42.785 ;
        RECT 128.465 42.615 128.635 42.785 ;
        RECT 128.925 42.615 129.095 42.785 ;
        RECT 129.385 42.615 129.555 42.785 ;
        RECT 129.845 42.615 130.015 42.785 ;
        RECT 130.305 42.615 130.475 42.785 ;
        RECT 130.765 42.615 130.935 42.785 ;
        RECT 131.225 42.615 131.395 42.785 ;
        RECT 131.685 42.615 131.855 42.785 ;
        RECT 132.145 42.615 132.315 42.785 ;
        RECT 132.605 42.615 132.775 42.785 ;
        RECT 133.065 42.615 133.235 42.785 ;
        RECT 133.525 42.615 133.695 42.785 ;
        RECT 133.985 42.615 134.155 42.785 ;
        RECT 134.445 42.615 134.615 42.785 ;
        RECT 134.905 42.615 135.075 42.785 ;
        RECT 135.365 42.615 135.535 42.785 ;
        RECT 135.825 42.615 135.995 42.785 ;
        RECT 136.285 42.615 136.455 42.785 ;
        RECT 136.745 42.615 136.915 42.785 ;
        RECT 137.205 42.615 137.375 42.785 ;
        RECT 137.665 42.615 137.835 42.785 ;
        RECT 138.125 42.615 138.295 42.785 ;
        RECT 138.585 42.615 138.755 42.785 ;
        RECT 139.045 42.615 139.215 42.785 ;
        RECT 139.505 42.615 139.675 42.785 ;
        RECT 139.965 42.615 140.135 42.785 ;
        RECT 140.425 42.615 140.595 42.785 ;
        RECT 140.885 42.615 141.055 42.785 ;
        RECT 141.345 42.615 141.515 42.785 ;
        RECT 141.805 42.615 141.975 42.785 ;
        RECT 142.265 42.615 142.435 42.785 ;
        RECT 142.725 42.615 142.895 42.785 ;
        RECT 143.185 42.615 143.355 42.785 ;
        RECT 143.645 42.615 143.815 42.785 ;
        RECT 144.105 42.615 144.275 42.785 ;
        RECT 144.565 42.615 144.735 42.785 ;
        RECT 145.025 42.615 145.195 42.785 ;
        RECT 145.485 42.615 145.655 42.785 ;
        RECT 145.945 42.615 146.115 42.785 ;
        RECT 146.405 42.615 146.575 42.785 ;
        RECT 146.865 42.615 147.035 42.785 ;
        RECT 147.325 42.615 147.495 42.785 ;
        RECT 147.785 42.615 147.955 42.785 ;
        RECT 148.245 42.615 148.415 42.785 ;
        RECT 148.705 42.615 148.875 42.785 ;
        RECT 149.165 42.615 149.335 42.785 ;
        RECT 149.625 42.615 149.795 42.785 ;
        RECT 150.085 42.615 150.255 42.785 ;
        RECT 150.545 42.615 150.715 42.785 ;
        RECT 151.005 42.615 151.175 42.785 ;
        RECT 151.465 42.615 151.635 42.785 ;
        RECT 151.925 42.615 152.095 42.785 ;
        RECT 92.585 41.085 92.755 41.255 ;
        RECT 93.505 40.405 93.675 40.575 ;
        RECT 99.025 41.085 99.195 41.255 ;
        RECT 100.405 41.425 100.575 41.595 ;
        RECT 139.045 42.105 139.215 42.275 ;
        RECT 139.045 41.085 139.215 41.255 ;
        RECT 139.965 41.085 140.135 41.255 ;
        RECT 141.345 41.085 141.515 41.255 ;
        RECT 141.810 41.085 141.980 41.255 ;
        RECT 142.215 41.765 142.385 41.935 ;
        RECT 142.725 41.425 142.895 41.595 ;
        RECT 144.105 41.765 144.275 41.935 ;
        RECT 143.645 41.085 143.815 41.255 ;
        RECT 147.225 41.765 147.395 41.935 ;
        RECT 145.365 40.745 145.535 40.915 ;
        RECT 147.225 41.085 147.395 41.255 ;
        RECT 148.305 41.060 148.475 41.230 ;
        RECT 148.605 40.745 148.775 40.915 ;
        RECT 150.085 40.405 150.255 40.575 ;
        RECT 91.205 39.895 91.375 40.065 ;
        RECT 91.665 39.895 91.835 40.065 ;
        RECT 92.125 39.895 92.295 40.065 ;
        RECT 92.585 39.895 92.755 40.065 ;
        RECT 93.045 39.895 93.215 40.065 ;
        RECT 93.505 39.895 93.675 40.065 ;
        RECT 93.965 39.895 94.135 40.065 ;
        RECT 94.425 39.895 94.595 40.065 ;
        RECT 94.885 39.895 95.055 40.065 ;
        RECT 95.345 39.895 95.515 40.065 ;
        RECT 95.805 39.895 95.975 40.065 ;
        RECT 96.265 39.895 96.435 40.065 ;
        RECT 96.725 39.895 96.895 40.065 ;
        RECT 97.185 39.895 97.355 40.065 ;
        RECT 97.645 39.895 97.815 40.065 ;
        RECT 98.105 39.895 98.275 40.065 ;
        RECT 98.565 39.895 98.735 40.065 ;
        RECT 99.025 39.895 99.195 40.065 ;
        RECT 99.485 39.895 99.655 40.065 ;
        RECT 99.945 39.895 100.115 40.065 ;
        RECT 100.405 39.895 100.575 40.065 ;
        RECT 100.865 39.895 101.035 40.065 ;
        RECT 101.325 39.895 101.495 40.065 ;
        RECT 101.785 39.895 101.955 40.065 ;
        RECT 102.245 39.895 102.415 40.065 ;
        RECT 102.705 39.895 102.875 40.065 ;
        RECT 103.165 39.895 103.335 40.065 ;
        RECT 103.625 39.895 103.795 40.065 ;
        RECT 104.085 39.895 104.255 40.065 ;
        RECT 104.545 39.895 104.715 40.065 ;
        RECT 105.005 39.895 105.175 40.065 ;
        RECT 105.465 39.895 105.635 40.065 ;
        RECT 105.925 39.895 106.095 40.065 ;
        RECT 106.385 39.895 106.555 40.065 ;
        RECT 106.845 39.895 107.015 40.065 ;
        RECT 107.305 39.895 107.475 40.065 ;
        RECT 107.765 39.895 107.935 40.065 ;
        RECT 108.225 39.895 108.395 40.065 ;
        RECT 108.685 39.895 108.855 40.065 ;
        RECT 109.145 39.895 109.315 40.065 ;
        RECT 109.605 39.895 109.775 40.065 ;
        RECT 110.065 39.895 110.235 40.065 ;
        RECT 110.525 39.895 110.695 40.065 ;
        RECT 110.985 39.895 111.155 40.065 ;
        RECT 111.445 39.895 111.615 40.065 ;
        RECT 111.905 39.895 112.075 40.065 ;
        RECT 112.365 39.895 112.535 40.065 ;
        RECT 112.825 39.895 112.995 40.065 ;
        RECT 113.285 39.895 113.455 40.065 ;
        RECT 113.745 39.895 113.915 40.065 ;
        RECT 114.205 39.895 114.375 40.065 ;
        RECT 114.665 39.895 114.835 40.065 ;
        RECT 115.125 39.895 115.295 40.065 ;
        RECT 115.585 39.895 115.755 40.065 ;
        RECT 116.045 39.895 116.215 40.065 ;
        RECT 116.505 39.895 116.675 40.065 ;
        RECT 116.965 39.895 117.135 40.065 ;
        RECT 117.425 39.895 117.595 40.065 ;
        RECT 117.885 39.895 118.055 40.065 ;
        RECT 118.345 39.895 118.515 40.065 ;
        RECT 118.805 39.895 118.975 40.065 ;
        RECT 119.265 39.895 119.435 40.065 ;
        RECT 119.725 39.895 119.895 40.065 ;
        RECT 120.185 39.895 120.355 40.065 ;
        RECT 120.645 39.895 120.815 40.065 ;
        RECT 121.105 39.895 121.275 40.065 ;
        RECT 121.565 39.895 121.735 40.065 ;
        RECT 122.025 39.895 122.195 40.065 ;
        RECT 122.485 39.895 122.655 40.065 ;
        RECT 122.945 39.895 123.115 40.065 ;
        RECT 123.405 39.895 123.575 40.065 ;
        RECT 123.865 39.895 124.035 40.065 ;
        RECT 124.325 39.895 124.495 40.065 ;
        RECT 124.785 39.895 124.955 40.065 ;
        RECT 125.245 39.895 125.415 40.065 ;
        RECT 125.705 39.895 125.875 40.065 ;
        RECT 126.165 39.895 126.335 40.065 ;
        RECT 126.625 39.895 126.795 40.065 ;
        RECT 127.085 39.895 127.255 40.065 ;
        RECT 127.545 39.895 127.715 40.065 ;
        RECT 128.005 39.895 128.175 40.065 ;
        RECT 128.465 39.895 128.635 40.065 ;
        RECT 128.925 39.895 129.095 40.065 ;
        RECT 129.385 39.895 129.555 40.065 ;
        RECT 129.845 39.895 130.015 40.065 ;
        RECT 130.305 39.895 130.475 40.065 ;
        RECT 130.765 39.895 130.935 40.065 ;
        RECT 131.225 39.895 131.395 40.065 ;
        RECT 131.685 39.895 131.855 40.065 ;
        RECT 132.145 39.895 132.315 40.065 ;
        RECT 132.605 39.895 132.775 40.065 ;
        RECT 133.065 39.895 133.235 40.065 ;
        RECT 133.525 39.895 133.695 40.065 ;
        RECT 133.985 39.895 134.155 40.065 ;
        RECT 134.445 39.895 134.615 40.065 ;
        RECT 134.905 39.895 135.075 40.065 ;
        RECT 135.365 39.895 135.535 40.065 ;
        RECT 135.825 39.895 135.995 40.065 ;
        RECT 136.285 39.895 136.455 40.065 ;
        RECT 136.745 39.895 136.915 40.065 ;
        RECT 137.205 39.895 137.375 40.065 ;
        RECT 137.665 39.895 137.835 40.065 ;
        RECT 138.125 39.895 138.295 40.065 ;
        RECT 138.585 39.895 138.755 40.065 ;
        RECT 139.045 39.895 139.215 40.065 ;
        RECT 139.505 39.895 139.675 40.065 ;
        RECT 139.965 39.895 140.135 40.065 ;
        RECT 140.425 39.895 140.595 40.065 ;
        RECT 140.885 39.895 141.055 40.065 ;
        RECT 141.345 39.895 141.515 40.065 ;
        RECT 141.805 39.895 141.975 40.065 ;
        RECT 142.265 39.895 142.435 40.065 ;
        RECT 142.725 39.895 142.895 40.065 ;
        RECT 143.185 39.895 143.355 40.065 ;
        RECT 143.645 39.895 143.815 40.065 ;
        RECT 144.105 39.895 144.275 40.065 ;
        RECT 144.565 39.895 144.735 40.065 ;
        RECT 145.025 39.895 145.195 40.065 ;
        RECT 145.485 39.895 145.655 40.065 ;
        RECT 145.945 39.895 146.115 40.065 ;
        RECT 146.405 39.895 146.575 40.065 ;
        RECT 146.865 39.895 147.035 40.065 ;
        RECT 147.325 39.895 147.495 40.065 ;
        RECT 147.785 39.895 147.955 40.065 ;
        RECT 148.245 39.895 148.415 40.065 ;
        RECT 148.705 39.895 148.875 40.065 ;
        RECT 149.165 39.895 149.335 40.065 ;
        RECT 149.625 39.895 149.795 40.065 ;
        RECT 150.085 39.895 150.255 40.065 ;
        RECT 150.545 39.895 150.715 40.065 ;
        RECT 151.005 39.895 151.175 40.065 ;
        RECT 151.465 39.895 151.635 40.065 ;
        RECT 151.925 39.895 152.095 40.065 ;
        RECT 6.055 37.350 6.275 37.570 ;
        RECT 102.245 39.385 102.415 39.555 ;
        RECT 99.945 38.705 100.115 38.875 ;
        RECT 98.565 38.025 98.735 38.195 ;
        RECT 99.025 37.685 99.195 37.855 ;
        RECT 101.325 37.685 101.495 37.855 ;
        RECT 106.385 39.385 106.555 39.555 ;
        RECT 108.225 38.705 108.395 38.875 ;
        RECT 109.605 38.705 109.775 38.875 ;
        RECT 110.065 38.705 110.235 38.875 ;
        RECT 105.925 38.025 106.095 38.195 ;
        RECT 110.985 38.705 111.155 38.875 ;
        RECT 108.685 37.685 108.855 37.855 ;
        RECT 111.905 38.025 112.075 38.195 ;
        RECT 111.445 37.685 111.615 37.855 ;
        RECT 113.745 39.045 113.915 39.215 ;
        RECT 114.665 38.365 114.835 38.535 ;
        RECT 115.585 38.365 115.755 38.535 ;
        RECT 115.125 37.685 115.295 37.855 ;
        RECT 119.265 38.365 119.435 38.535 ;
        RECT 120.185 38.705 120.355 38.875 ;
        RECT 120.645 38.025 120.815 38.195 ;
        RECT 121.565 38.705 121.735 38.875 ;
        RECT 122.485 38.705 122.655 38.875 ;
        RECT 123.405 38.705 123.575 38.875 ;
        RECT 123.865 39.045 124.035 39.215 ;
        RECT 124.325 38.705 124.495 38.875 ;
        RECT 121.105 38.025 121.275 38.195 ;
        RECT 125.705 38.705 125.875 38.875 ;
        RECT 126.625 38.705 126.795 38.875 ;
        RECT 127.085 38.705 127.255 38.875 ;
        RECT 127.545 38.705 127.715 38.875 ;
        RECT 125.245 38.025 125.415 38.195 ;
        RECT 128.925 38.705 129.095 38.875 ;
        RECT 129.845 38.705 130.015 38.875 ;
        RECT 128.465 37.685 128.635 37.855 ;
        RECT 129.845 37.685 130.015 37.855 ;
        RECT 136.745 39.385 136.915 39.555 ;
        RECT 132.605 38.705 132.775 38.875 ;
        RECT 131.225 38.025 131.395 38.195 ;
        RECT 132.145 37.685 132.315 37.855 ;
        RECT 140.425 39.385 140.595 39.555 ;
        RECT 137.495 38.705 137.665 38.875 ;
        RECT 139.045 38.365 139.215 38.535 ;
        RECT 139.965 38.705 140.135 38.875 ;
        RECT 139.505 38.365 139.675 38.535 ;
        RECT 141.345 39.045 141.515 39.215 ;
        RECT 141.345 38.025 141.515 38.195 ;
        RECT 144.105 38.705 144.275 38.875 ;
        RECT 143.645 38.365 143.815 38.535 ;
        RECT 147.325 38.705 147.495 38.875 ;
        RECT 145.945 37.685 146.115 37.855 ;
        RECT 150.085 38.705 150.255 38.875 ;
        RECT 91.205 37.175 91.375 37.345 ;
        RECT 91.665 37.175 91.835 37.345 ;
        RECT 92.125 37.175 92.295 37.345 ;
        RECT 92.585 37.175 92.755 37.345 ;
        RECT 93.045 37.175 93.215 37.345 ;
        RECT 93.505 37.175 93.675 37.345 ;
        RECT 93.965 37.175 94.135 37.345 ;
        RECT 94.425 37.175 94.595 37.345 ;
        RECT 94.885 37.175 95.055 37.345 ;
        RECT 95.345 37.175 95.515 37.345 ;
        RECT 95.805 37.175 95.975 37.345 ;
        RECT 96.265 37.175 96.435 37.345 ;
        RECT 96.725 37.175 96.895 37.345 ;
        RECT 97.185 37.175 97.355 37.345 ;
        RECT 97.645 37.175 97.815 37.345 ;
        RECT 98.105 37.175 98.275 37.345 ;
        RECT 98.565 37.175 98.735 37.345 ;
        RECT 99.025 37.175 99.195 37.345 ;
        RECT 99.485 37.175 99.655 37.345 ;
        RECT 99.945 37.175 100.115 37.345 ;
        RECT 100.405 37.175 100.575 37.345 ;
        RECT 100.865 37.175 101.035 37.345 ;
        RECT 101.325 37.175 101.495 37.345 ;
        RECT 101.785 37.175 101.955 37.345 ;
        RECT 102.245 37.175 102.415 37.345 ;
        RECT 102.705 37.175 102.875 37.345 ;
        RECT 103.165 37.175 103.335 37.345 ;
        RECT 103.625 37.175 103.795 37.345 ;
        RECT 104.085 37.175 104.255 37.345 ;
        RECT 104.545 37.175 104.715 37.345 ;
        RECT 105.005 37.175 105.175 37.345 ;
        RECT 105.465 37.175 105.635 37.345 ;
        RECT 105.925 37.175 106.095 37.345 ;
        RECT 106.385 37.175 106.555 37.345 ;
        RECT 106.845 37.175 107.015 37.345 ;
        RECT 107.305 37.175 107.475 37.345 ;
        RECT 107.765 37.175 107.935 37.345 ;
        RECT 108.225 37.175 108.395 37.345 ;
        RECT 108.685 37.175 108.855 37.345 ;
        RECT 109.145 37.175 109.315 37.345 ;
        RECT 109.605 37.175 109.775 37.345 ;
        RECT 110.065 37.175 110.235 37.345 ;
        RECT 110.525 37.175 110.695 37.345 ;
        RECT 110.985 37.175 111.155 37.345 ;
        RECT 111.445 37.175 111.615 37.345 ;
        RECT 111.905 37.175 112.075 37.345 ;
        RECT 112.365 37.175 112.535 37.345 ;
        RECT 112.825 37.175 112.995 37.345 ;
        RECT 113.285 37.175 113.455 37.345 ;
        RECT 113.745 37.175 113.915 37.345 ;
        RECT 114.205 37.175 114.375 37.345 ;
        RECT 114.665 37.175 114.835 37.345 ;
        RECT 115.125 37.175 115.295 37.345 ;
        RECT 115.585 37.175 115.755 37.345 ;
        RECT 116.045 37.175 116.215 37.345 ;
        RECT 116.505 37.175 116.675 37.345 ;
        RECT 116.965 37.175 117.135 37.345 ;
        RECT 117.425 37.175 117.595 37.345 ;
        RECT 117.885 37.175 118.055 37.345 ;
        RECT 118.345 37.175 118.515 37.345 ;
        RECT 118.805 37.175 118.975 37.345 ;
        RECT 119.265 37.175 119.435 37.345 ;
        RECT 119.725 37.175 119.895 37.345 ;
        RECT 120.185 37.175 120.355 37.345 ;
        RECT 120.645 37.175 120.815 37.345 ;
        RECT 121.105 37.175 121.275 37.345 ;
        RECT 121.565 37.175 121.735 37.345 ;
        RECT 122.025 37.175 122.195 37.345 ;
        RECT 122.485 37.175 122.655 37.345 ;
        RECT 122.945 37.175 123.115 37.345 ;
        RECT 123.405 37.175 123.575 37.345 ;
        RECT 123.865 37.175 124.035 37.345 ;
        RECT 124.325 37.175 124.495 37.345 ;
        RECT 124.785 37.175 124.955 37.345 ;
        RECT 125.245 37.175 125.415 37.345 ;
        RECT 125.705 37.175 125.875 37.345 ;
        RECT 126.165 37.175 126.335 37.345 ;
        RECT 126.625 37.175 126.795 37.345 ;
        RECT 127.085 37.175 127.255 37.345 ;
        RECT 127.545 37.175 127.715 37.345 ;
        RECT 128.005 37.175 128.175 37.345 ;
        RECT 128.465 37.175 128.635 37.345 ;
        RECT 128.925 37.175 129.095 37.345 ;
        RECT 129.385 37.175 129.555 37.345 ;
        RECT 129.845 37.175 130.015 37.345 ;
        RECT 130.305 37.175 130.475 37.345 ;
        RECT 130.765 37.175 130.935 37.345 ;
        RECT 131.225 37.175 131.395 37.345 ;
        RECT 131.685 37.175 131.855 37.345 ;
        RECT 132.145 37.175 132.315 37.345 ;
        RECT 132.605 37.175 132.775 37.345 ;
        RECT 133.065 37.175 133.235 37.345 ;
        RECT 133.525 37.175 133.695 37.345 ;
        RECT 133.985 37.175 134.155 37.345 ;
        RECT 134.445 37.175 134.615 37.345 ;
        RECT 134.905 37.175 135.075 37.345 ;
        RECT 135.365 37.175 135.535 37.345 ;
        RECT 135.825 37.175 135.995 37.345 ;
        RECT 136.285 37.175 136.455 37.345 ;
        RECT 136.745 37.175 136.915 37.345 ;
        RECT 137.205 37.175 137.375 37.345 ;
        RECT 137.665 37.175 137.835 37.345 ;
        RECT 138.125 37.175 138.295 37.345 ;
        RECT 138.585 37.175 138.755 37.345 ;
        RECT 139.045 37.175 139.215 37.345 ;
        RECT 139.505 37.175 139.675 37.345 ;
        RECT 139.965 37.175 140.135 37.345 ;
        RECT 140.425 37.175 140.595 37.345 ;
        RECT 140.885 37.175 141.055 37.345 ;
        RECT 141.345 37.175 141.515 37.345 ;
        RECT 141.805 37.175 141.975 37.345 ;
        RECT 142.265 37.175 142.435 37.345 ;
        RECT 142.725 37.175 142.895 37.345 ;
        RECT 143.185 37.175 143.355 37.345 ;
        RECT 143.645 37.175 143.815 37.345 ;
        RECT 144.105 37.175 144.275 37.345 ;
        RECT 144.565 37.175 144.735 37.345 ;
        RECT 145.025 37.175 145.195 37.345 ;
        RECT 145.485 37.175 145.655 37.345 ;
        RECT 145.945 37.175 146.115 37.345 ;
        RECT 146.405 37.175 146.575 37.345 ;
        RECT 146.865 37.175 147.035 37.345 ;
        RECT 147.325 37.175 147.495 37.345 ;
        RECT 147.785 37.175 147.955 37.345 ;
        RECT 148.245 37.175 148.415 37.345 ;
        RECT 148.705 37.175 148.875 37.345 ;
        RECT 149.165 37.175 149.335 37.345 ;
        RECT 149.625 37.175 149.795 37.345 ;
        RECT 150.085 37.175 150.255 37.345 ;
        RECT 150.545 37.175 150.715 37.345 ;
        RECT 151.005 37.175 151.175 37.345 ;
        RECT 151.465 37.175 151.635 37.345 ;
        RECT 151.925 37.175 152.095 37.345 ;
        RECT 93.965 36.665 94.135 36.835 ;
        RECT 92.585 35.645 92.755 35.815 ;
        RECT 95.345 36.325 95.515 36.495 ;
        RECT 97.185 36.665 97.355 36.835 ;
        RECT 98.105 36.325 98.275 36.495 ;
        RECT 99.025 36.665 99.195 36.835 ;
        RECT 94.885 34.965 95.055 35.135 ;
        RECT 98.565 35.645 98.735 35.815 ;
        RECT 97.185 34.965 97.355 35.135 ;
        RECT 99.945 34.965 100.115 35.135 ;
        RECT 100.405 35.305 100.575 35.475 ;
        RECT 100.865 35.645 101.035 35.815 ;
        RECT 103.165 36.325 103.335 36.495 ;
        RECT 102.705 35.645 102.875 35.815 ;
        RECT 102.245 34.965 102.415 35.135 ;
        RECT 104.545 35.645 104.715 35.815 ;
        RECT 105.925 35.985 106.095 36.155 ;
        RECT 108.225 36.665 108.395 36.835 ;
        RECT 105.465 35.645 105.635 35.815 ;
        RECT 107.305 35.645 107.475 35.815 ;
        RECT 109.605 35.645 109.775 35.815 ;
        RECT 113.285 36.665 113.455 36.835 ;
        RECT 110.525 35.645 110.695 35.815 ;
        RECT 110.985 35.645 111.155 35.815 ;
        RECT 112.365 35.645 112.535 35.815 ;
        RECT 114.205 35.985 114.375 36.155 ;
        RECT 115.125 36.325 115.295 36.495 ;
        RECT 114.665 35.645 114.835 35.815 ;
        RECT 117.425 35.985 117.595 36.155 ;
        RECT 120.645 36.665 120.815 36.835 ;
        RECT 116.045 35.645 116.215 35.815 ;
        RECT 117.885 35.645 118.055 35.815 ;
        RECT 122.485 36.665 122.655 36.835 ;
        RECT 121.105 35.985 121.275 36.155 ;
        RECT 121.565 35.645 121.735 35.815 ;
        RECT 120.185 35.305 120.355 35.475 ;
        RECT 123.570 35.645 123.740 35.815 ;
        RECT 122.945 34.965 123.115 35.135 ;
        RECT 125.705 35.985 125.875 36.155 ;
        RECT 126.165 35.645 126.335 35.815 ;
        RECT 130.305 36.665 130.475 36.835 ;
        RECT 127.545 35.645 127.715 35.815 ;
        RECT 128.005 35.305 128.175 35.475 ;
        RECT 128.465 35.645 128.635 35.815 ;
        RECT 129.385 35.645 129.555 35.815 ;
        RECT 126.625 34.965 126.795 35.135 ;
        RECT 132.605 36.325 132.775 36.495 ;
        RECT 136.745 36.665 136.915 36.835 ;
        RECT 131.225 35.645 131.395 35.815 ;
        RECT 132.975 35.645 133.145 35.815 ;
        RECT 133.525 35.645 133.695 35.815 ;
        RECT 133.990 35.645 134.160 35.815 ;
        RECT 134.905 35.305 135.075 35.475 ;
        RECT 135.365 35.645 135.535 35.815 ;
        RECT 135.850 35.645 136.020 35.815 ;
        RECT 138.125 35.985 138.295 36.155 ;
        RECT 140.425 36.665 140.595 36.835 ;
        RECT 137.665 35.645 137.835 35.815 ;
        RECT 138.585 35.645 138.755 35.815 ;
        RECT 139.965 35.645 140.135 35.815 ;
        RECT 141.345 35.985 141.515 36.155 ;
        RECT 141.810 35.645 141.980 35.815 ;
        RECT 142.215 36.325 142.385 36.495 ;
        RECT 142.725 35.305 142.895 35.475 ;
        RECT 144.105 36.325 144.275 36.495 ;
        RECT 143.645 35.645 143.815 35.815 ;
        RECT 147.225 36.325 147.395 36.495 ;
        RECT 145.365 35.305 145.535 35.475 ;
        RECT 147.225 35.645 147.395 35.815 ;
        RECT 150.085 36.665 150.255 36.835 ;
        RECT 148.305 35.620 148.475 35.790 ;
        RECT 148.605 35.305 148.775 35.475 ;
        RECT 6.110 32.025 6.300 34.010 ;
        RECT 59.135 32.590 59.325 34.575 ;
        RECT 91.205 34.455 91.375 34.625 ;
        RECT 91.665 34.455 91.835 34.625 ;
        RECT 92.125 34.455 92.295 34.625 ;
        RECT 92.585 34.455 92.755 34.625 ;
        RECT 93.045 34.455 93.215 34.625 ;
        RECT 93.505 34.455 93.675 34.625 ;
        RECT 93.965 34.455 94.135 34.625 ;
        RECT 94.425 34.455 94.595 34.625 ;
        RECT 94.885 34.455 95.055 34.625 ;
        RECT 95.345 34.455 95.515 34.625 ;
        RECT 95.805 34.455 95.975 34.625 ;
        RECT 96.265 34.455 96.435 34.625 ;
        RECT 96.725 34.455 96.895 34.625 ;
        RECT 97.185 34.455 97.355 34.625 ;
        RECT 97.645 34.455 97.815 34.625 ;
        RECT 98.105 34.455 98.275 34.625 ;
        RECT 98.565 34.455 98.735 34.625 ;
        RECT 99.025 34.455 99.195 34.625 ;
        RECT 99.485 34.455 99.655 34.625 ;
        RECT 99.945 34.455 100.115 34.625 ;
        RECT 100.405 34.455 100.575 34.625 ;
        RECT 100.865 34.455 101.035 34.625 ;
        RECT 101.325 34.455 101.495 34.625 ;
        RECT 101.785 34.455 101.955 34.625 ;
        RECT 102.245 34.455 102.415 34.625 ;
        RECT 102.705 34.455 102.875 34.625 ;
        RECT 103.165 34.455 103.335 34.625 ;
        RECT 103.625 34.455 103.795 34.625 ;
        RECT 104.085 34.455 104.255 34.625 ;
        RECT 104.545 34.455 104.715 34.625 ;
        RECT 105.005 34.455 105.175 34.625 ;
        RECT 105.465 34.455 105.635 34.625 ;
        RECT 105.925 34.455 106.095 34.625 ;
        RECT 106.385 34.455 106.555 34.625 ;
        RECT 106.845 34.455 107.015 34.625 ;
        RECT 107.305 34.455 107.475 34.625 ;
        RECT 107.765 34.455 107.935 34.625 ;
        RECT 108.225 34.455 108.395 34.625 ;
        RECT 108.685 34.455 108.855 34.625 ;
        RECT 109.145 34.455 109.315 34.625 ;
        RECT 109.605 34.455 109.775 34.625 ;
        RECT 110.065 34.455 110.235 34.625 ;
        RECT 110.525 34.455 110.695 34.625 ;
        RECT 110.985 34.455 111.155 34.625 ;
        RECT 111.445 34.455 111.615 34.625 ;
        RECT 111.905 34.455 112.075 34.625 ;
        RECT 112.365 34.455 112.535 34.625 ;
        RECT 112.825 34.455 112.995 34.625 ;
        RECT 113.285 34.455 113.455 34.625 ;
        RECT 113.745 34.455 113.915 34.625 ;
        RECT 114.205 34.455 114.375 34.625 ;
        RECT 114.665 34.455 114.835 34.625 ;
        RECT 115.125 34.455 115.295 34.625 ;
        RECT 115.585 34.455 115.755 34.625 ;
        RECT 116.045 34.455 116.215 34.625 ;
        RECT 116.505 34.455 116.675 34.625 ;
        RECT 116.965 34.455 117.135 34.625 ;
        RECT 117.425 34.455 117.595 34.625 ;
        RECT 117.885 34.455 118.055 34.625 ;
        RECT 118.345 34.455 118.515 34.625 ;
        RECT 118.805 34.455 118.975 34.625 ;
        RECT 119.265 34.455 119.435 34.625 ;
        RECT 119.725 34.455 119.895 34.625 ;
        RECT 120.185 34.455 120.355 34.625 ;
        RECT 120.645 34.455 120.815 34.625 ;
        RECT 121.105 34.455 121.275 34.625 ;
        RECT 121.565 34.455 121.735 34.625 ;
        RECT 122.025 34.455 122.195 34.625 ;
        RECT 122.485 34.455 122.655 34.625 ;
        RECT 122.945 34.455 123.115 34.625 ;
        RECT 123.405 34.455 123.575 34.625 ;
        RECT 123.865 34.455 124.035 34.625 ;
        RECT 124.325 34.455 124.495 34.625 ;
        RECT 124.785 34.455 124.955 34.625 ;
        RECT 125.245 34.455 125.415 34.625 ;
        RECT 125.705 34.455 125.875 34.625 ;
        RECT 126.165 34.455 126.335 34.625 ;
        RECT 126.625 34.455 126.795 34.625 ;
        RECT 127.085 34.455 127.255 34.625 ;
        RECT 127.545 34.455 127.715 34.625 ;
        RECT 128.005 34.455 128.175 34.625 ;
        RECT 128.465 34.455 128.635 34.625 ;
        RECT 128.925 34.455 129.095 34.625 ;
        RECT 129.385 34.455 129.555 34.625 ;
        RECT 129.845 34.455 130.015 34.625 ;
        RECT 130.305 34.455 130.475 34.625 ;
        RECT 130.765 34.455 130.935 34.625 ;
        RECT 131.225 34.455 131.395 34.625 ;
        RECT 131.685 34.455 131.855 34.625 ;
        RECT 132.145 34.455 132.315 34.625 ;
        RECT 132.605 34.455 132.775 34.625 ;
        RECT 133.065 34.455 133.235 34.625 ;
        RECT 133.525 34.455 133.695 34.625 ;
        RECT 133.985 34.455 134.155 34.625 ;
        RECT 134.445 34.455 134.615 34.625 ;
        RECT 134.905 34.455 135.075 34.625 ;
        RECT 135.365 34.455 135.535 34.625 ;
        RECT 135.825 34.455 135.995 34.625 ;
        RECT 136.285 34.455 136.455 34.625 ;
        RECT 136.745 34.455 136.915 34.625 ;
        RECT 137.205 34.455 137.375 34.625 ;
        RECT 137.665 34.455 137.835 34.625 ;
        RECT 138.125 34.455 138.295 34.625 ;
        RECT 138.585 34.455 138.755 34.625 ;
        RECT 139.045 34.455 139.215 34.625 ;
        RECT 139.505 34.455 139.675 34.625 ;
        RECT 139.965 34.455 140.135 34.625 ;
        RECT 140.425 34.455 140.595 34.625 ;
        RECT 140.885 34.455 141.055 34.625 ;
        RECT 141.345 34.455 141.515 34.625 ;
        RECT 141.805 34.455 141.975 34.625 ;
        RECT 142.265 34.455 142.435 34.625 ;
        RECT 142.725 34.455 142.895 34.625 ;
        RECT 143.185 34.455 143.355 34.625 ;
        RECT 143.645 34.455 143.815 34.625 ;
        RECT 144.105 34.455 144.275 34.625 ;
        RECT 144.565 34.455 144.735 34.625 ;
        RECT 145.025 34.455 145.195 34.625 ;
        RECT 145.485 34.455 145.655 34.625 ;
        RECT 145.945 34.455 146.115 34.625 ;
        RECT 146.405 34.455 146.575 34.625 ;
        RECT 146.865 34.455 147.035 34.625 ;
        RECT 147.325 34.455 147.495 34.625 ;
        RECT 147.785 34.455 147.955 34.625 ;
        RECT 148.245 34.455 148.415 34.625 ;
        RECT 148.705 34.455 148.875 34.625 ;
        RECT 149.165 34.455 149.335 34.625 ;
        RECT 149.625 34.455 149.795 34.625 ;
        RECT 150.085 34.455 150.255 34.625 ;
        RECT 150.545 34.455 150.715 34.625 ;
        RECT 151.005 34.455 151.175 34.625 ;
        RECT 151.465 34.455 151.635 34.625 ;
        RECT 151.925 34.455 152.095 34.625 ;
        RECT 100.405 33.945 100.575 34.115 ;
        RECT 98.105 33.265 98.275 33.435 ;
        RECT 99.485 32.245 99.655 32.415 ;
        RECT 100.865 33.945 101.035 34.115 ;
        RECT 103.165 33.265 103.335 33.435 ;
        RECT 102.705 32.245 102.875 32.415 ;
        RECT 105.465 33.605 105.635 33.775 ;
        RECT 104.925 33.295 105.095 33.465 ;
        RECT 107.765 33.945 107.935 34.115 ;
        RECT 105.925 33.265 106.095 33.435 ;
        RECT 106.845 33.265 107.015 33.435 ;
        RECT 107.305 33.265 107.475 33.435 ;
        RECT 104.085 32.245 104.255 32.415 ;
        RECT 108.225 32.585 108.395 32.755 ;
        RECT 111.905 33.605 112.075 33.775 ;
        RECT 110.065 33.265 110.235 33.435 ;
        RECT 110.985 33.265 111.155 33.435 ;
        RECT 112.365 33.265 112.535 33.435 ;
        RECT 112.825 33.265 112.995 33.435 ;
        RECT 114.205 32.925 114.375 33.095 ;
        RECT 115.125 33.265 115.295 33.435 ;
        RECT 116.045 33.605 116.215 33.775 ;
        RECT 120.185 33.945 120.355 34.115 ;
        RECT 117.885 33.265 118.055 33.435 ;
        RECT 119.265 33.265 119.435 33.435 ;
        RECT 118.805 32.925 118.975 33.095 ;
        RECT 122.025 33.945 122.195 34.115 ;
        RECT 123.405 33.605 123.575 33.775 ;
        RECT 125.245 33.945 125.415 34.115 ;
        RECT 122.485 33.265 122.655 33.435 ;
        RECT 122.945 33.265 123.115 33.435 ;
        RECT 124.325 33.265 124.495 33.435 ;
        RECT 117.885 32.245 118.055 32.415 ;
        RECT 127.545 33.605 127.715 33.775 ;
        RECT 126.625 33.265 126.795 33.435 ;
        RECT 128.005 33.265 128.175 33.435 ;
        RECT 128.465 33.265 128.635 33.435 ;
        RECT 133.985 33.945 134.155 34.115 ;
        RECT 131.225 33.265 131.395 33.435 ;
        RECT 132.605 33.265 132.775 33.435 ;
        RECT 133.065 33.265 133.235 33.435 ;
        RECT 131.685 32.585 131.855 32.755 ;
        RECT 146.865 33.945 147.035 34.115 ;
        RECT 146.405 33.265 146.575 33.435 ;
        RECT 148.245 33.945 148.415 34.115 ;
        RECT 147.325 33.265 147.495 33.435 ;
        RECT 147.785 33.265 147.955 33.435 ;
        RECT 150.545 33.265 150.715 33.435 ;
        RECT 149.625 32.585 149.795 32.755 ;
        RECT 91.205 31.735 91.375 31.905 ;
        RECT 91.665 31.735 91.835 31.905 ;
        RECT 92.125 31.735 92.295 31.905 ;
        RECT 92.585 31.735 92.755 31.905 ;
        RECT 93.045 31.735 93.215 31.905 ;
        RECT 93.505 31.735 93.675 31.905 ;
        RECT 93.965 31.735 94.135 31.905 ;
        RECT 94.425 31.735 94.595 31.905 ;
        RECT 94.885 31.735 95.055 31.905 ;
        RECT 95.345 31.735 95.515 31.905 ;
        RECT 95.805 31.735 95.975 31.905 ;
        RECT 96.265 31.735 96.435 31.905 ;
        RECT 96.725 31.735 96.895 31.905 ;
        RECT 97.185 31.735 97.355 31.905 ;
        RECT 97.645 31.735 97.815 31.905 ;
        RECT 98.105 31.735 98.275 31.905 ;
        RECT 98.565 31.735 98.735 31.905 ;
        RECT 99.025 31.735 99.195 31.905 ;
        RECT 99.485 31.735 99.655 31.905 ;
        RECT 99.945 31.735 100.115 31.905 ;
        RECT 100.405 31.735 100.575 31.905 ;
        RECT 100.865 31.735 101.035 31.905 ;
        RECT 101.325 31.735 101.495 31.905 ;
        RECT 101.785 31.735 101.955 31.905 ;
        RECT 102.245 31.735 102.415 31.905 ;
        RECT 102.705 31.735 102.875 31.905 ;
        RECT 103.165 31.735 103.335 31.905 ;
        RECT 103.625 31.735 103.795 31.905 ;
        RECT 104.085 31.735 104.255 31.905 ;
        RECT 104.545 31.735 104.715 31.905 ;
        RECT 105.005 31.735 105.175 31.905 ;
        RECT 105.465 31.735 105.635 31.905 ;
        RECT 105.925 31.735 106.095 31.905 ;
        RECT 106.385 31.735 106.555 31.905 ;
        RECT 106.845 31.735 107.015 31.905 ;
        RECT 107.305 31.735 107.475 31.905 ;
        RECT 107.765 31.735 107.935 31.905 ;
        RECT 108.225 31.735 108.395 31.905 ;
        RECT 108.685 31.735 108.855 31.905 ;
        RECT 109.145 31.735 109.315 31.905 ;
        RECT 109.605 31.735 109.775 31.905 ;
        RECT 110.065 31.735 110.235 31.905 ;
        RECT 110.525 31.735 110.695 31.905 ;
        RECT 110.985 31.735 111.155 31.905 ;
        RECT 111.445 31.735 111.615 31.905 ;
        RECT 111.905 31.735 112.075 31.905 ;
        RECT 112.365 31.735 112.535 31.905 ;
        RECT 112.825 31.735 112.995 31.905 ;
        RECT 113.285 31.735 113.455 31.905 ;
        RECT 113.745 31.735 113.915 31.905 ;
        RECT 114.205 31.735 114.375 31.905 ;
        RECT 114.665 31.735 114.835 31.905 ;
        RECT 115.125 31.735 115.295 31.905 ;
        RECT 115.585 31.735 115.755 31.905 ;
        RECT 116.045 31.735 116.215 31.905 ;
        RECT 116.505 31.735 116.675 31.905 ;
        RECT 116.965 31.735 117.135 31.905 ;
        RECT 117.425 31.735 117.595 31.905 ;
        RECT 117.885 31.735 118.055 31.905 ;
        RECT 118.345 31.735 118.515 31.905 ;
        RECT 118.805 31.735 118.975 31.905 ;
        RECT 119.265 31.735 119.435 31.905 ;
        RECT 119.725 31.735 119.895 31.905 ;
        RECT 120.185 31.735 120.355 31.905 ;
        RECT 120.645 31.735 120.815 31.905 ;
        RECT 121.105 31.735 121.275 31.905 ;
        RECT 121.565 31.735 121.735 31.905 ;
        RECT 122.025 31.735 122.195 31.905 ;
        RECT 122.485 31.735 122.655 31.905 ;
        RECT 122.945 31.735 123.115 31.905 ;
        RECT 123.405 31.735 123.575 31.905 ;
        RECT 123.865 31.735 124.035 31.905 ;
        RECT 124.325 31.735 124.495 31.905 ;
        RECT 124.785 31.735 124.955 31.905 ;
        RECT 125.245 31.735 125.415 31.905 ;
        RECT 125.705 31.735 125.875 31.905 ;
        RECT 126.165 31.735 126.335 31.905 ;
        RECT 126.625 31.735 126.795 31.905 ;
        RECT 127.085 31.735 127.255 31.905 ;
        RECT 127.545 31.735 127.715 31.905 ;
        RECT 128.005 31.735 128.175 31.905 ;
        RECT 128.465 31.735 128.635 31.905 ;
        RECT 128.925 31.735 129.095 31.905 ;
        RECT 129.385 31.735 129.555 31.905 ;
        RECT 129.845 31.735 130.015 31.905 ;
        RECT 130.305 31.735 130.475 31.905 ;
        RECT 130.765 31.735 130.935 31.905 ;
        RECT 131.225 31.735 131.395 31.905 ;
        RECT 131.685 31.735 131.855 31.905 ;
        RECT 132.145 31.735 132.315 31.905 ;
        RECT 132.605 31.735 132.775 31.905 ;
        RECT 133.065 31.735 133.235 31.905 ;
        RECT 133.525 31.735 133.695 31.905 ;
        RECT 133.985 31.735 134.155 31.905 ;
        RECT 134.445 31.735 134.615 31.905 ;
        RECT 134.905 31.735 135.075 31.905 ;
        RECT 135.365 31.735 135.535 31.905 ;
        RECT 135.825 31.735 135.995 31.905 ;
        RECT 136.285 31.735 136.455 31.905 ;
        RECT 136.745 31.735 136.915 31.905 ;
        RECT 137.205 31.735 137.375 31.905 ;
        RECT 137.665 31.735 137.835 31.905 ;
        RECT 138.125 31.735 138.295 31.905 ;
        RECT 138.585 31.735 138.755 31.905 ;
        RECT 139.045 31.735 139.215 31.905 ;
        RECT 139.505 31.735 139.675 31.905 ;
        RECT 139.965 31.735 140.135 31.905 ;
        RECT 140.425 31.735 140.595 31.905 ;
        RECT 140.885 31.735 141.055 31.905 ;
        RECT 141.345 31.735 141.515 31.905 ;
        RECT 141.805 31.735 141.975 31.905 ;
        RECT 142.265 31.735 142.435 31.905 ;
        RECT 142.725 31.735 142.895 31.905 ;
        RECT 143.185 31.735 143.355 31.905 ;
        RECT 143.645 31.735 143.815 31.905 ;
        RECT 144.105 31.735 144.275 31.905 ;
        RECT 144.565 31.735 144.735 31.905 ;
        RECT 145.025 31.735 145.195 31.905 ;
        RECT 145.485 31.735 145.655 31.905 ;
        RECT 145.945 31.735 146.115 31.905 ;
        RECT 146.405 31.735 146.575 31.905 ;
        RECT 146.865 31.735 147.035 31.905 ;
        RECT 147.325 31.735 147.495 31.905 ;
        RECT 147.785 31.735 147.955 31.905 ;
        RECT 148.245 31.735 148.415 31.905 ;
        RECT 148.705 31.735 148.875 31.905 ;
        RECT 149.165 31.735 149.335 31.905 ;
        RECT 149.625 31.735 149.795 31.905 ;
        RECT 150.085 31.735 150.255 31.905 ;
        RECT 150.545 31.735 150.715 31.905 ;
        RECT 151.005 31.735 151.175 31.905 ;
        RECT 151.465 31.735 151.635 31.905 ;
        RECT 151.925 31.735 152.095 31.905 ;
        RECT 6.110 28.870 6.300 30.855 ;
        RECT 93.505 31.225 93.675 31.395 ;
        RECT 92.585 30.205 92.755 30.375 ;
        RECT 8.050 28.940 8.415 29.470 ;
        RECT 99.485 31.225 99.655 31.395 ;
        RECT 98.565 30.205 98.735 30.375 ;
        RECT 107.305 31.225 107.475 31.395 ;
        RECT 106.385 30.205 106.555 30.375 ;
        RECT 115.125 31.225 115.295 31.395 ;
        RECT 114.205 30.205 114.375 30.375 ;
        RECT 119.265 30.205 119.435 30.375 ;
        RECT 119.725 30.205 119.895 30.375 ;
        RECT 122.025 30.885 122.195 31.055 ;
        RECT 122.945 30.205 123.115 30.375 ;
        RECT 130.305 31.225 130.475 31.395 ;
        RECT 131.225 30.205 131.395 30.375 ;
        RECT 137.665 31.225 137.835 31.395 ;
        RECT 138.585 30.205 138.755 30.375 ;
        RECT 143.185 30.205 143.355 30.375 ;
        RECT 144.565 30.545 144.735 30.715 ;
        RECT 149.625 31.225 149.795 31.395 ;
        RECT 150.085 29.865 150.255 30.035 ;
        RECT 91.205 29.015 91.375 29.185 ;
        RECT 91.665 29.015 91.835 29.185 ;
        RECT 92.125 29.015 92.295 29.185 ;
        RECT 92.585 29.015 92.755 29.185 ;
        RECT 93.045 29.015 93.215 29.185 ;
        RECT 93.505 29.015 93.675 29.185 ;
        RECT 93.965 29.015 94.135 29.185 ;
        RECT 94.425 29.015 94.595 29.185 ;
        RECT 94.885 29.015 95.055 29.185 ;
        RECT 95.345 29.015 95.515 29.185 ;
        RECT 95.805 29.015 95.975 29.185 ;
        RECT 96.265 29.015 96.435 29.185 ;
        RECT 96.725 29.015 96.895 29.185 ;
        RECT 97.185 29.015 97.355 29.185 ;
        RECT 97.645 29.015 97.815 29.185 ;
        RECT 98.105 29.015 98.275 29.185 ;
        RECT 98.565 29.015 98.735 29.185 ;
        RECT 99.025 29.015 99.195 29.185 ;
        RECT 99.485 29.015 99.655 29.185 ;
        RECT 99.945 29.015 100.115 29.185 ;
        RECT 100.405 29.015 100.575 29.185 ;
        RECT 100.865 29.015 101.035 29.185 ;
        RECT 101.325 29.015 101.495 29.185 ;
        RECT 101.785 29.015 101.955 29.185 ;
        RECT 102.245 29.015 102.415 29.185 ;
        RECT 102.705 29.015 102.875 29.185 ;
        RECT 103.165 29.015 103.335 29.185 ;
        RECT 103.625 29.015 103.795 29.185 ;
        RECT 104.085 29.015 104.255 29.185 ;
        RECT 104.545 29.015 104.715 29.185 ;
        RECT 105.005 29.015 105.175 29.185 ;
        RECT 105.465 29.015 105.635 29.185 ;
        RECT 105.925 29.015 106.095 29.185 ;
        RECT 106.385 29.015 106.555 29.185 ;
        RECT 106.845 29.015 107.015 29.185 ;
        RECT 107.305 29.015 107.475 29.185 ;
        RECT 107.765 29.015 107.935 29.185 ;
        RECT 108.225 29.015 108.395 29.185 ;
        RECT 108.685 29.015 108.855 29.185 ;
        RECT 109.145 29.015 109.315 29.185 ;
        RECT 109.605 29.015 109.775 29.185 ;
        RECT 110.065 29.015 110.235 29.185 ;
        RECT 110.525 29.015 110.695 29.185 ;
        RECT 110.985 29.015 111.155 29.185 ;
        RECT 111.445 29.015 111.615 29.185 ;
        RECT 111.905 29.015 112.075 29.185 ;
        RECT 112.365 29.015 112.535 29.185 ;
        RECT 112.825 29.015 112.995 29.185 ;
        RECT 113.285 29.015 113.455 29.185 ;
        RECT 113.745 29.015 113.915 29.185 ;
        RECT 114.205 29.015 114.375 29.185 ;
        RECT 114.665 29.015 114.835 29.185 ;
        RECT 115.125 29.015 115.295 29.185 ;
        RECT 115.585 29.015 115.755 29.185 ;
        RECT 116.045 29.015 116.215 29.185 ;
        RECT 116.505 29.015 116.675 29.185 ;
        RECT 116.965 29.015 117.135 29.185 ;
        RECT 117.425 29.015 117.595 29.185 ;
        RECT 117.885 29.015 118.055 29.185 ;
        RECT 118.345 29.015 118.515 29.185 ;
        RECT 118.805 29.015 118.975 29.185 ;
        RECT 119.265 29.015 119.435 29.185 ;
        RECT 119.725 29.015 119.895 29.185 ;
        RECT 120.185 29.015 120.355 29.185 ;
        RECT 120.645 29.015 120.815 29.185 ;
        RECT 121.105 29.015 121.275 29.185 ;
        RECT 121.565 29.015 121.735 29.185 ;
        RECT 122.025 29.015 122.195 29.185 ;
        RECT 122.485 29.015 122.655 29.185 ;
        RECT 122.945 29.015 123.115 29.185 ;
        RECT 123.405 29.015 123.575 29.185 ;
        RECT 123.865 29.015 124.035 29.185 ;
        RECT 124.325 29.015 124.495 29.185 ;
        RECT 124.785 29.015 124.955 29.185 ;
        RECT 125.245 29.015 125.415 29.185 ;
        RECT 125.705 29.015 125.875 29.185 ;
        RECT 126.165 29.015 126.335 29.185 ;
        RECT 126.625 29.015 126.795 29.185 ;
        RECT 127.085 29.015 127.255 29.185 ;
        RECT 127.545 29.015 127.715 29.185 ;
        RECT 128.005 29.015 128.175 29.185 ;
        RECT 128.465 29.015 128.635 29.185 ;
        RECT 128.925 29.015 129.095 29.185 ;
        RECT 129.385 29.015 129.555 29.185 ;
        RECT 129.845 29.015 130.015 29.185 ;
        RECT 130.305 29.015 130.475 29.185 ;
        RECT 130.765 29.015 130.935 29.185 ;
        RECT 131.225 29.015 131.395 29.185 ;
        RECT 131.685 29.015 131.855 29.185 ;
        RECT 132.145 29.015 132.315 29.185 ;
        RECT 132.605 29.015 132.775 29.185 ;
        RECT 133.065 29.015 133.235 29.185 ;
        RECT 133.525 29.015 133.695 29.185 ;
        RECT 133.985 29.015 134.155 29.185 ;
        RECT 134.445 29.015 134.615 29.185 ;
        RECT 134.905 29.015 135.075 29.185 ;
        RECT 135.365 29.015 135.535 29.185 ;
        RECT 135.825 29.015 135.995 29.185 ;
        RECT 136.285 29.015 136.455 29.185 ;
        RECT 136.745 29.015 136.915 29.185 ;
        RECT 137.205 29.015 137.375 29.185 ;
        RECT 137.665 29.015 137.835 29.185 ;
        RECT 138.125 29.015 138.295 29.185 ;
        RECT 138.585 29.015 138.755 29.185 ;
        RECT 139.045 29.015 139.215 29.185 ;
        RECT 139.505 29.015 139.675 29.185 ;
        RECT 139.965 29.015 140.135 29.185 ;
        RECT 140.425 29.015 140.595 29.185 ;
        RECT 140.885 29.015 141.055 29.185 ;
        RECT 141.345 29.015 141.515 29.185 ;
        RECT 141.805 29.015 141.975 29.185 ;
        RECT 142.265 29.015 142.435 29.185 ;
        RECT 142.725 29.015 142.895 29.185 ;
        RECT 143.185 29.015 143.355 29.185 ;
        RECT 143.645 29.015 143.815 29.185 ;
        RECT 144.105 29.015 144.275 29.185 ;
        RECT 144.565 29.015 144.735 29.185 ;
        RECT 145.025 29.015 145.195 29.185 ;
        RECT 145.485 29.015 145.655 29.185 ;
        RECT 145.945 29.015 146.115 29.185 ;
        RECT 146.405 29.015 146.575 29.185 ;
        RECT 146.865 29.015 147.035 29.185 ;
        RECT 147.325 29.015 147.495 29.185 ;
        RECT 147.785 29.015 147.955 29.185 ;
        RECT 148.245 29.015 148.415 29.185 ;
        RECT 148.705 29.015 148.875 29.185 ;
        RECT 149.165 29.015 149.335 29.185 ;
        RECT 149.625 29.015 149.795 29.185 ;
        RECT 150.085 29.015 150.255 29.185 ;
        RECT 150.545 29.015 150.715 29.185 ;
        RECT 151.005 29.015 151.175 29.185 ;
        RECT 151.465 29.015 151.635 29.185 ;
        RECT 151.925 29.015 152.095 29.185 ;
        RECT 6.100 19.865 6.290 21.850 ;
        RECT 59.135 24.435 59.325 26.420 ;
        RECT 59.095 20.600 59.375 20.880 ;
        RECT 6.100 16.710 6.290 18.695 ;
        RECT 8.560 16.620 9.610 17.985 ;
        RECT 59.140 10.515 59.330 12.500 ;
        RECT 53.335 8.005 53.805 8.460 ;
        RECT 59.140 7.860 59.330 9.845 ;
      LAYER met1 ;
        RECT 84.840 222.455 85.360 222.940 ;
        RECT 88.500 222.470 89.020 222.955 ;
        RECT 85.005 200.565 85.160 222.455 ;
        RECT 84.920 200.305 85.240 200.565 ;
        RECT 1.005 194.685 2.505 195.185 ;
        RECT 1.005 194.670 69.085 194.685 ;
        RECT 1.005 194.190 119.550 194.670 ;
        RECT 1.005 194.185 69.410 194.190 ;
        RECT 1.005 193.685 2.505 194.185 ;
        RECT 68.930 189.230 69.410 194.185 ;
        RECT 80.520 193.990 80.840 194.050 ;
        RECT 81.915 193.990 82.205 194.035 ;
        RECT 80.520 193.850 82.205 193.990 ;
        RECT 80.520 193.790 80.840 193.850 ;
        RECT 81.915 193.805 82.205 193.850 ;
        RECT 110.420 193.990 110.740 194.050 ;
        RECT 111.815 193.990 112.105 194.035 ;
        RECT 110.420 193.850 112.105 193.990 ;
        RECT 110.420 193.790 110.740 193.850 ;
        RECT 111.815 193.805 112.105 193.850 ;
        RECT 86.960 192.970 87.280 193.030 ;
        RECT 88.815 192.970 89.105 193.015 ;
        RECT 86.960 192.830 89.105 192.970 ;
        RECT 86.960 192.770 87.280 192.830 ;
        RECT 88.815 192.785 89.105 192.830 ;
        RECT 81.440 192.430 81.760 192.690 ;
        RECT 100.300 192.430 100.620 192.690 ;
        RECT 101.235 192.630 101.525 192.675 ;
        RECT 102.600 192.630 102.920 192.690 ;
        RECT 101.235 192.490 102.920 192.630 ;
        RECT 101.235 192.445 101.525 192.490 ;
        RECT 102.600 192.430 102.920 192.490 ;
        RECT 111.340 192.430 111.660 192.690 ;
        RECT 82.360 192.290 82.680 192.350 ;
        RECT 86.055 192.290 86.345 192.335 ;
        RECT 82.360 192.150 86.345 192.290 ;
        RECT 82.360 192.090 82.680 192.150 ;
        RECT 86.055 192.105 86.345 192.150 ;
        RECT 102.155 192.290 102.445 192.335 ;
        RECT 106.740 192.290 107.060 192.350 ;
        RECT 102.155 192.150 107.060 192.290 ;
        RECT 102.155 192.105 102.445 192.150 ;
        RECT 106.740 192.090 107.060 192.150 ;
        RECT 71.250 191.470 121.935 191.950 ;
        RECT 77.315 191.270 77.605 191.315 ;
        RECT 81.440 191.270 81.760 191.330 ;
        RECT 106.280 191.270 106.600 191.330 ;
        RECT 77.315 191.130 81.760 191.270 ;
        RECT 77.315 191.085 77.605 191.130 ;
        RECT 81.440 191.070 81.760 191.130 ;
        RECT 95.330 191.130 106.600 191.270 ;
        RECT 92.650 190.930 92.940 190.975 ;
        RECT 94.335 190.930 94.625 190.975 ;
        RECT 92.650 190.790 94.625 190.930 ;
        RECT 92.650 190.745 92.940 190.790 ;
        RECT 94.335 190.745 94.625 190.790 ;
        RECT 70.400 190.590 70.720 190.650 ;
        RECT 72.715 190.590 73.005 190.635 ;
        RECT 70.400 190.450 73.005 190.590 ;
        RECT 70.400 190.390 70.720 190.450 ;
        RECT 72.715 190.405 73.005 190.450 ;
        RECT 80.980 190.390 81.300 190.650 ;
        RECT 82.820 190.390 83.140 190.650 ;
        RECT 95.330 190.635 95.470 191.130 ;
        RECT 106.280 191.070 106.600 191.130 ;
        RECT 110.895 191.270 111.185 191.315 ;
        RECT 111.340 191.270 111.660 191.330 ;
        RECT 110.895 191.130 111.660 191.270 ;
        RECT 110.895 191.085 111.185 191.130 ;
        RECT 111.340 191.070 111.660 191.130 ;
        RECT 107.660 190.930 107.980 190.990 ;
        RECT 95.790 190.790 107.980 190.930 ;
        RECT 95.790 190.635 95.930 190.790 ;
        RECT 107.660 190.730 107.980 190.790 ;
        RECT 83.755 190.590 84.045 190.635 ;
        RECT 83.755 190.450 94.550 190.590 ;
        RECT 83.755 190.405 84.045 190.450 ;
        RECT 79.570 190.250 79.860 190.295 ;
        RECT 81.910 190.250 82.200 190.295 ;
        RECT 79.570 190.110 82.200 190.250 ;
        RECT 79.570 190.065 79.860 190.110 ;
        RECT 81.910 190.065 82.200 190.110 ;
        RECT 82.375 190.250 82.665 190.295 ;
        RECT 87.880 190.250 88.200 190.310 ;
        RECT 94.410 190.295 94.550 190.450 ;
        RECT 95.255 190.405 95.545 190.635 ;
        RECT 95.715 190.405 96.005 190.635 ;
        RECT 100.300 190.590 100.620 190.650 ;
        RECT 102.155 190.590 102.445 190.635 ;
        RECT 100.300 190.450 102.445 190.590 ;
        RECT 100.300 190.390 100.620 190.450 ;
        RECT 102.155 190.405 102.445 190.450 ;
        RECT 103.060 190.390 103.380 190.650 ;
        RECT 103.535 190.590 103.825 190.635 ;
        RECT 104.440 190.590 104.760 190.650 ;
        RECT 103.535 190.450 104.760 190.590 ;
        RECT 103.535 190.405 103.825 190.450 ;
        RECT 104.440 190.390 104.760 190.450 ;
        RECT 105.835 190.405 106.125 190.635 ;
        RECT 107.215 190.590 107.505 190.635 ;
        RECT 109.040 190.590 109.360 190.650 ;
        RECT 107.215 190.450 109.360 190.590 ;
        RECT 107.215 190.405 107.505 190.450 ;
        RECT 82.375 190.110 88.200 190.250 ;
        RECT 82.375 190.065 82.665 190.110 ;
        RECT 87.880 190.050 88.200 190.110 ;
        RECT 89.285 190.250 89.575 190.295 ;
        RECT 91.805 190.250 92.095 190.295 ;
        RECT 92.995 190.250 93.285 190.295 ;
        RECT 89.285 190.110 93.285 190.250 ;
        RECT 89.285 190.065 89.575 190.110 ;
        RECT 91.805 190.065 92.095 190.110 ;
        RECT 92.995 190.065 93.285 190.110 ;
        RECT 93.875 190.065 94.165 190.295 ;
        RECT 94.335 190.065 94.625 190.295 ;
        RECT 94.780 190.250 95.100 190.310 ;
        RECT 100.775 190.250 101.065 190.295 ;
        RECT 103.980 190.250 104.300 190.310 ;
        RECT 94.780 190.110 104.300 190.250 ;
        RECT 80.075 189.910 80.365 189.955 ;
        RECT 81.450 189.910 81.740 189.955 ;
        RECT 80.075 189.770 81.740 189.910 ;
        RECT 80.075 189.725 80.365 189.770 ;
        RECT 81.450 189.725 81.740 189.770 ;
        RECT 83.740 189.910 84.060 189.970 ;
        RECT 89.720 189.910 90.010 189.955 ;
        RECT 91.290 189.910 91.580 189.955 ;
        RECT 93.390 189.910 93.680 189.955 ;
        RECT 83.740 189.770 89.490 189.910 ;
        RECT 83.740 189.710 84.060 189.770 ;
        RECT 73.620 189.370 73.940 189.630 ;
        RECT 83.295 189.570 83.585 189.615 ;
        RECT 84.200 189.570 84.520 189.630 ;
        RECT 83.295 189.430 84.520 189.570 ;
        RECT 83.295 189.385 83.585 189.430 ;
        RECT 84.200 189.370 84.520 189.430 ;
        RECT 86.960 189.370 87.280 189.630 ;
        RECT 89.350 189.570 89.490 189.770 ;
        RECT 89.720 189.770 93.680 189.910 ;
        RECT 89.720 189.725 90.010 189.770 ;
        RECT 91.290 189.725 91.580 189.770 ;
        RECT 93.390 189.725 93.680 189.770 ;
        RECT 93.950 189.630 94.090 190.065 ;
        RECT 94.410 189.910 94.550 190.065 ;
        RECT 94.780 190.050 95.100 190.110 ;
        RECT 100.775 190.065 101.065 190.110 ;
        RECT 103.980 190.050 104.300 190.110 ;
        RECT 101.235 189.910 101.525 189.955 ;
        RECT 94.410 189.770 101.525 189.910 ;
        RECT 101.235 189.725 101.525 189.770 ;
        RECT 93.860 189.570 94.180 189.630 ;
        RECT 89.350 189.430 94.180 189.570 ;
        RECT 93.860 189.370 94.180 189.430 ;
        RECT 94.320 189.570 94.640 189.630 ;
        RECT 97.555 189.570 97.845 189.615 ;
        RECT 94.320 189.430 97.845 189.570 ;
        RECT 94.320 189.370 94.640 189.430 ;
        RECT 97.555 189.385 97.845 189.430 ;
        RECT 103.520 189.570 103.840 189.630 ;
        RECT 105.910 189.570 106.050 190.405 ;
        RECT 109.040 190.390 109.360 190.450 ;
        RECT 117.795 190.590 118.085 190.635 ;
        RECT 117.795 190.450 120.310 190.590 ;
        RECT 117.795 190.405 118.085 190.450 ;
        RECT 106.300 190.250 106.590 190.295 ;
        RECT 108.640 190.250 108.930 190.295 ;
        RECT 106.300 190.110 108.930 190.250 ;
        RECT 106.300 190.065 106.590 190.110 ;
        RECT 108.640 190.065 108.930 190.110 ;
        RECT 120.170 189.970 120.310 190.450 ;
        RECT 106.760 189.910 107.050 189.955 ;
        RECT 108.135 189.910 108.425 189.955 ;
        RECT 106.760 189.770 108.425 189.910 ;
        RECT 106.760 189.725 107.050 189.770 ;
        RECT 108.135 189.725 108.425 189.770 ;
        RECT 120.080 189.710 120.400 189.970 ;
        RECT 103.520 189.430 106.050 189.570 ;
        RECT 111.800 189.570 112.120 189.630 ;
        RECT 116.875 189.570 117.165 189.615 ;
        RECT 111.800 189.430 117.165 189.570 ;
        RECT 103.520 189.370 103.840 189.430 ;
        RECT 111.800 189.370 112.120 189.430 ;
        RECT 116.875 189.385 117.165 189.430 ;
        RECT 68.930 188.750 119.550 189.230 ;
        RECT 68.930 183.790 69.410 188.750 ;
        RECT 73.620 188.350 73.940 188.610 ;
        RECT 82.360 188.350 82.680 188.610 ;
        RECT 82.820 188.550 83.140 188.610 ;
        RECT 83.755 188.550 84.045 188.595 ;
        RECT 94.320 188.550 94.640 188.610 ;
        RECT 82.820 188.410 84.045 188.550 ;
        RECT 82.820 188.350 83.140 188.410 ;
        RECT 83.755 188.365 84.045 188.410 ;
        RECT 84.750 188.410 94.640 188.550 ;
        RECT 73.710 187.530 73.850 188.350 ;
        RECT 84.750 188.210 84.890 188.410 ;
        RECT 94.320 188.350 94.640 188.410 ;
        RECT 103.980 188.350 104.300 188.610 ;
        RECT 107.660 188.350 107.980 188.610 ;
        RECT 112.735 188.550 113.025 188.595 ;
        RECT 119.160 188.550 119.480 188.610 ;
        RECT 112.735 188.410 119.480 188.550 ;
        RECT 112.735 188.365 113.025 188.410 ;
        RECT 82.450 188.070 84.890 188.210 ;
        RECT 85.160 188.210 85.450 188.255 ;
        RECT 87.260 188.210 87.550 188.255 ;
        RECT 88.830 188.210 89.120 188.255 ;
        RECT 85.160 188.070 89.120 188.210 ;
        RECT 82.450 187.915 82.590 188.070 ;
        RECT 85.160 188.025 85.450 188.070 ;
        RECT 87.260 188.025 87.550 188.070 ;
        RECT 88.830 188.025 89.120 188.070 ;
        RECT 97.580 188.210 97.870 188.255 ;
        RECT 99.680 188.210 99.970 188.255 ;
        RECT 101.250 188.210 101.540 188.255 ;
        RECT 97.580 188.070 101.540 188.210 ;
        RECT 97.580 188.025 97.870 188.070 ;
        RECT 99.680 188.025 99.970 188.070 ;
        RECT 101.250 188.025 101.540 188.070 ;
        RECT 106.280 188.010 106.600 188.270 ;
        RECT 82.375 187.685 82.665 187.915 ;
        RECT 84.675 187.685 84.965 187.915 ;
        RECT 85.555 187.870 85.845 187.915 ;
        RECT 86.745 187.870 87.035 187.915 ;
        RECT 89.265 187.870 89.555 187.915 ;
        RECT 85.555 187.730 89.555 187.870 ;
        RECT 85.555 187.685 85.845 187.730 ;
        RECT 86.745 187.685 87.035 187.730 ;
        RECT 89.265 187.685 89.555 187.730 ;
        RECT 93.860 187.870 94.180 187.930 ;
        RECT 97.095 187.870 97.385 187.915 ;
        RECT 93.860 187.730 97.385 187.870 ;
        RECT 80.535 187.530 80.825 187.575 ;
        RECT 73.710 187.390 80.825 187.530 ;
        RECT 80.535 187.345 80.825 187.390 ;
        RECT 82.820 187.540 83.110 187.575 ;
        RECT 82.820 187.400 83.510 187.540 ;
        RECT 82.820 187.345 83.110 187.400 ;
        RECT 83.370 186.850 83.510 187.400 ;
        RECT 83.740 187.530 84.060 187.590 ;
        RECT 84.750 187.530 84.890 187.685 ;
        RECT 93.860 187.670 94.180 187.730 ;
        RECT 97.095 187.685 97.385 187.730 ;
        RECT 97.975 187.870 98.265 187.915 ;
        RECT 99.165 187.870 99.455 187.915 ;
        RECT 101.685 187.870 101.975 187.915 ;
        RECT 97.975 187.730 101.975 187.870 ;
        RECT 97.975 187.685 98.265 187.730 ;
        RECT 99.165 187.685 99.455 187.730 ;
        RECT 101.685 187.685 101.975 187.730 ;
        RECT 104.440 187.670 104.760 187.930 ;
        RECT 105.835 187.870 106.125 187.915 ;
        RECT 108.120 187.870 108.440 187.930 ;
        RECT 111.800 187.870 112.120 187.930 ;
        RECT 105.835 187.730 112.120 187.870 ;
        RECT 105.835 187.685 106.125 187.730 ;
        RECT 83.740 187.390 84.890 187.530 ;
        RECT 83.740 187.330 84.060 187.390 ;
        RECT 94.780 187.330 95.100 187.590 ;
        RECT 95.715 187.530 96.005 187.575 ;
        RECT 99.840 187.530 100.160 187.590 ;
        RECT 104.530 187.530 104.670 187.670 ;
        RECT 95.715 187.390 104.670 187.530 ;
        RECT 95.715 187.345 96.005 187.390 ;
        RECT 84.200 187.190 84.520 187.250 ;
        RECT 85.900 187.190 86.190 187.235 ;
        RECT 84.200 187.050 86.190 187.190 ;
        RECT 84.200 186.990 84.520 187.050 ;
        RECT 85.900 187.005 86.190 187.050 ;
        RECT 89.260 187.190 89.580 187.250 ;
        RECT 92.035 187.190 92.325 187.235 ;
        RECT 89.260 187.050 92.325 187.190 ;
        RECT 89.260 186.990 89.580 187.050 ;
        RECT 92.035 187.005 92.325 187.050 ;
        RECT 85.120 186.850 85.440 186.910 ;
        RECT 91.575 186.850 91.865 186.895 ;
        RECT 95.790 186.850 95.930 187.345 ;
        RECT 99.840 187.330 100.160 187.390 ;
        RECT 105.375 187.345 105.665 187.575 ;
        RECT 98.460 187.235 98.780 187.250 ;
        RECT 98.430 187.005 98.780 187.235 ;
        RECT 98.460 186.990 98.780 187.005 ;
        RECT 101.220 187.190 101.540 187.250 ;
        RECT 104.455 187.190 104.745 187.235 ;
        RECT 101.220 187.050 104.745 187.190 ;
        RECT 105.450 187.190 105.590 187.345 ;
        RECT 106.740 187.330 107.060 187.590 ;
        RECT 107.750 187.575 107.890 187.730 ;
        RECT 108.120 187.670 108.440 187.730 ;
        RECT 111.800 187.670 112.120 187.730 ;
        RECT 107.675 187.345 107.965 187.575 ;
        RECT 108.595 187.345 108.885 187.575 ;
        RECT 111.355 187.530 111.645 187.575 ;
        RECT 111.890 187.530 112.030 187.670 ;
        RECT 111.355 187.390 112.030 187.530 ;
        RECT 111.355 187.345 111.645 187.390 ;
        RECT 108.670 187.190 108.810 187.345 ;
        RECT 112.810 187.190 112.950 188.365 ;
        RECT 119.160 188.350 119.480 188.410 ;
        RECT 113.655 187.870 113.945 187.915 ;
        RECT 113.655 187.730 115.250 187.870 ;
        RECT 113.655 187.685 113.945 187.730 ;
        RECT 115.110 187.575 115.250 187.730 ;
        RECT 115.035 187.345 115.325 187.575 ;
        RECT 105.450 187.050 112.950 187.190 ;
        RECT 101.220 186.990 101.540 187.050 ;
        RECT 104.455 187.005 104.745 187.050 ;
        RECT 83.370 186.710 95.930 186.850 ;
        RECT 96.175 186.850 96.465 186.895 ;
        RECT 102.600 186.850 102.920 186.910 ;
        RECT 96.175 186.710 102.920 186.850 ;
        RECT 85.120 186.650 85.440 186.710 ;
        RECT 91.575 186.665 91.865 186.710 ;
        RECT 96.175 186.665 96.465 186.710 ;
        RECT 102.600 186.650 102.920 186.710 ;
        RECT 113.180 186.850 113.500 186.910 ;
        RECT 114.115 186.850 114.405 186.895 ;
        RECT 113.180 186.710 114.405 186.850 ;
        RECT 113.180 186.650 113.500 186.710 ;
        RECT 114.115 186.665 114.405 186.710 ;
        RECT 121.455 186.510 121.935 191.470 ;
        RECT 71.250 186.030 121.935 186.510 ;
        RECT 79.140 185.830 79.460 185.890 ;
        RECT 83.740 185.830 84.060 185.890 ;
        RECT 79.140 185.690 84.060 185.830 ;
        RECT 79.140 185.630 79.460 185.690 ;
        RECT 83.740 185.630 84.060 185.690 ;
        RECT 89.260 185.630 89.580 185.890 ;
        RECT 98.460 185.630 98.780 185.890 ;
        RECT 98.920 185.830 99.240 185.890 ;
        RECT 99.395 185.830 99.685 185.875 ;
        RECT 103.520 185.830 103.840 185.890 ;
        RECT 98.920 185.690 103.840 185.830 ;
        RECT 98.920 185.630 99.240 185.690 ;
        RECT 99.395 185.645 99.685 185.690 ;
        RECT 103.520 185.630 103.840 185.690 ;
        RECT 103.995 185.830 104.285 185.875 ;
        RECT 106.280 185.830 106.600 185.890 ;
        RECT 103.995 185.690 106.600 185.830 ;
        RECT 103.995 185.645 104.285 185.690 ;
        RECT 106.280 185.630 106.600 185.690 ;
        RECT 108.120 185.630 108.440 185.890 ;
        RECT 85.120 184.950 85.440 185.210 ;
        RECT 86.515 185.150 86.805 185.195 ;
        RECT 89.350 185.150 89.490 185.630 ;
        RECT 94.410 185.350 102.370 185.490 ;
        RECT 94.410 185.210 94.550 185.350 ;
        RECT 86.515 185.010 89.490 185.150 ;
        RECT 86.515 184.965 86.805 185.010 ;
        RECT 94.320 184.950 94.640 185.210 ;
        RECT 99.380 185.150 99.670 185.195 ;
        RECT 101.220 185.150 101.540 185.210 ;
        RECT 102.230 185.195 102.370 185.350 ;
        RECT 99.380 185.010 101.540 185.150 ;
        RECT 99.380 184.965 99.670 185.010 ;
        RECT 101.220 184.950 101.540 185.010 ;
        RECT 102.155 184.965 102.445 185.195 ;
        RECT 102.600 184.950 102.920 185.210 ;
        RECT 103.060 184.950 103.380 185.210 ;
        RECT 107.215 185.150 107.505 185.195 ;
        RECT 108.210 185.150 108.350 185.630 ;
        RECT 112.230 185.490 112.520 185.535 ;
        RECT 113.180 185.490 113.500 185.550 ;
        RECT 112.230 185.350 113.500 185.490 ;
        RECT 112.230 185.305 112.520 185.350 ;
        RECT 113.180 185.290 113.500 185.350 ;
        RECT 108.595 185.150 108.885 185.195 ;
        RECT 107.215 185.010 107.890 185.150 ;
        RECT 108.210 185.010 108.885 185.150 ;
        RECT 107.215 184.965 107.505 185.010 ;
        RECT 87.880 184.810 88.200 184.870 ;
        RECT 89.735 184.810 90.025 184.855 ;
        RECT 87.880 184.670 90.025 184.810 ;
        RECT 87.880 184.610 88.200 184.670 ;
        RECT 89.735 184.625 90.025 184.670 ;
        RECT 91.100 184.610 91.420 184.870 ;
        RECT 93.875 184.810 94.165 184.855 ;
        RECT 100.300 184.810 100.620 184.870 ;
        RECT 93.875 184.670 100.620 184.810 ;
        RECT 93.875 184.625 94.165 184.670 ;
        RECT 100.300 184.610 100.620 184.670 ;
        RECT 101.695 184.810 101.985 184.855 ;
        RECT 103.150 184.810 103.290 184.950 ;
        RECT 101.695 184.670 103.290 184.810 ;
        RECT 101.695 184.625 101.985 184.670 ;
        RECT 106.280 184.610 106.600 184.870 ;
        RECT 86.960 184.470 87.280 184.530 ;
        RECT 92.940 184.470 93.260 184.530 ;
        RECT 101.235 184.470 101.525 184.515 ;
        RECT 106.370 184.470 106.510 184.610 ;
        RECT 107.750 184.515 107.890 185.010 ;
        RECT 108.595 184.965 108.885 185.010 ;
        RECT 110.880 184.610 111.200 184.870 ;
        RECT 111.775 184.810 112.065 184.855 ;
        RECT 112.965 184.810 113.255 184.855 ;
        RECT 115.485 184.810 115.775 184.855 ;
        RECT 111.775 184.670 115.775 184.810 ;
        RECT 111.775 184.625 112.065 184.670 ;
        RECT 112.965 184.625 113.255 184.670 ;
        RECT 115.485 184.625 115.775 184.670 ;
        RECT 86.130 184.330 97.310 184.470 ;
        RECT 83.740 183.930 84.060 184.190 ;
        RECT 86.130 184.175 86.270 184.330 ;
        RECT 86.960 184.270 87.280 184.330 ;
        RECT 92.940 184.270 93.260 184.330 ;
        RECT 86.055 183.945 86.345 184.175 ;
        RECT 95.700 184.130 96.020 184.190 ;
        RECT 96.635 184.130 96.925 184.175 ;
        RECT 95.700 183.990 96.925 184.130 ;
        RECT 97.170 184.130 97.310 184.330 ;
        RECT 101.235 184.330 106.510 184.470 ;
        RECT 101.235 184.285 101.525 184.330 ;
        RECT 107.675 184.285 107.965 184.515 ;
        RECT 111.380 184.470 111.670 184.515 ;
        RECT 113.480 184.470 113.770 184.515 ;
        RECT 115.050 184.470 115.340 184.515 ;
        RECT 111.380 184.330 115.340 184.470 ;
        RECT 111.380 184.285 111.670 184.330 ;
        RECT 113.480 184.285 113.770 184.330 ;
        RECT 115.050 184.285 115.340 184.330 ;
        RECT 102.155 184.130 102.445 184.175 ;
        RECT 97.170 183.990 102.445 184.130 ;
        RECT 95.700 183.930 96.020 183.990 ;
        RECT 96.635 183.945 96.925 183.990 ;
        RECT 102.155 183.945 102.445 183.990 ;
        RECT 106.295 184.130 106.585 184.175 ;
        RECT 106.740 184.130 107.060 184.190 ;
        RECT 106.295 183.990 107.060 184.130 ;
        RECT 106.295 183.945 106.585 183.990 ;
        RECT 106.740 183.930 107.060 183.990 ;
        RECT 117.795 184.130 118.085 184.175 ;
        RECT 117.795 183.990 119.850 184.130 ;
        RECT 117.795 183.945 118.085 183.990 ;
        RECT 68.930 183.310 119.550 183.790 ;
        RECT 68.930 178.350 69.410 183.310 ;
        RECT 83.740 182.910 84.060 183.170 ;
        RECT 87.880 182.910 88.200 183.170 ;
        RECT 90.195 183.110 90.485 183.155 ;
        RECT 91.100 183.110 91.420 183.170 ;
        RECT 90.195 182.970 91.420 183.110 ;
        RECT 90.195 182.925 90.485 182.970 ;
        RECT 91.100 182.910 91.420 182.970 ;
        RECT 93.875 183.110 94.165 183.155 ;
        RECT 94.320 183.110 94.640 183.170 ;
        RECT 93.875 182.970 94.640 183.110 ;
        RECT 93.875 182.925 94.165 182.970 ;
        RECT 94.320 182.910 94.640 182.970 ;
        RECT 83.830 182.430 83.970 182.910 ;
        RECT 87.970 182.770 88.110 182.910 ;
        RECT 98.920 182.770 99.240 182.830 ;
        RECT 87.970 182.630 99.240 182.770 ;
        RECT 86.975 182.430 87.265 182.475 ;
        RECT 83.830 182.290 87.265 182.430 ;
        RECT 86.975 182.245 87.265 182.290 ;
        RECT 92.495 182.090 92.785 182.135 ;
        RECT 92.940 182.090 93.260 182.150 ;
        RECT 92.495 181.950 93.260 182.090 ;
        RECT 92.495 181.905 92.785 181.950 ;
        RECT 92.940 181.890 93.260 181.950 ;
        RECT 95.700 181.890 96.020 182.150 ;
        RECT 96.710 182.135 96.850 182.630 ;
        RECT 98.920 182.570 99.240 182.630 ;
        RECT 117.795 182.430 118.085 182.475 ;
        RECT 119.710 182.430 119.850 183.990 ;
        RECT 117.795 182.290 119.850 182.430 ;
        RECT 117.795 182.245 118.085 182.290 ;
        RECT 96.635 181.905 96.925 182.135 ;
        RECT 114.115 182.090 114.405 182.135 ;
        RECT 114.575 182.090 114.865 182.135 ;
        RECT 114.115 181.950 114.865 182.090 ;
        RECT 114.115 181.905 114.405 181.950 ;
        RECT 114.575 181.905 114.865 181.950 ;
        RECT 93.860 181.750 94.180 181.810 ;
        RECT 97.555 181.750 97.845 181.795 ;
        RECT 93.860 181.610 97.845 181.750 ;
        RECT 93.860 181.550 94.180 181.610 ;
        RECT 97.555 181.565 97.845 181.610 ;
        RECT 102.600 181.750 102.920 181.810 ;
        RECT 103.995 181.750 104.285 181.795 ;
        RECT 102.600 181.610 104.285 181.750 ;
        RECT 102.600 181.550 102.920 181.610 ;
        RECT 103.995 181.565 104.285 181.610 ;
        RECT 104.915 181.565 105.205 181.795 ;
        RECT 105.820 181.750 106.140 181.810 ;
        RECT 115.020 181.750 115.340 181.810 ;
        RECT 105.820 181.610 115.340 181.750 ;
        RECT 94.795 181.410 95.085 181.455 ;
        RECT 100.300 181.410 100.620 181.470 ;
        RECT 94.795 181.270 100.620 181.410 ;
        RECT 104.990 181.410 105.130 181.565 ;
        RECT 105.820 181.550 106.140 181.610 ;
        RECT 115.020 181.550 115.340 181.610 ;
        RECT 106.280 181.410 106.600 181.470 ;
        RECT 104.990 181.270 106.600 181.410 ;
        RECT 94.795 181.225 95.085 181.270 ;
        RECT 100.300 181.210 100.620 181.270 ;
        RECT 106.280 181.210 106.600 181.270 ;
        RECT 111.800 181.410 112.120 181.470 ;
        RECT 113.655 181.410 113.945 181.455 ;
        RECT 111.800 181.270 113.945 181.410 ;
        RECT 111.800 181.210 112.120 181.270 ;
        RECT 113.655 181.225 113.945 181.270 ;
        RECT 121.455 181.070 121.935 186.030 ;
        RECT 71.250 180.590 121.935 181.070 ;
        RECT 99.380 180.390 99.700 180.450 ;
        RECT 98.550 180.250 99.700 180.390 ;
        RECT 98.550 180.095 98.690 180.250 ;
        RECT 99.380 180.190 99.700 180.250 ;
        RECT 101.235 180.390 101.525 180.435 ;
        RECT 107.660 180.390 107.980 180.450 ;
        RECT 101.235 180.250 107.980 180.390 ;
        RECT 101.235 180.205 101.525 180.250 ;
        RECT 107.660 180.190 107.980 180.250 ;
        RECT 110.880 180.190 111.200 180.450 ;
        RECT 77.295 180.050 77.945 180.095 ;
        RECT 80.895 180.050 81.185 180.095 ;
        RECT 77.295 179.910 81.185 180.050 ;
        RECT 77.295 179.865 77.945 179.910 ;
        RECT 80.595 179.865 81.185 179.910 ;
        RECT 98.475 179.865 98.765 180.095 ;
        RECT 99.840 180.050 100.160 180.110 ;
        RECT 110.970 180.050 111.110 180.190 ;
        RECT 99.840 179.910 111.110 180.050 ;
        RECT 73.620 179.510 73.940 179.770 ;
        RECT 74.100 179.710 74.390 179.755 ;
        RECT 75.935 179.710 76.225 179.755 ;
        RECT 79.515 179.710 79.805 179.755 ;
        RECT 74.100 179.570 79.805 179.710 ;
        RECT 74.100 179.525 74.390 179.570 ;
        RECT 75.935 179.525 76.225 179.570 ;
        RECT 79.515 179.525 79.805 179.570 ;
        RECT 80.595 179.710 80.885 179.865 ;
        RECT 82.360 179.710 82.680 179.770 ;
        RECT 86.055 179.710 86.345 179.755 ;
        RECT 80.595 179.570 82.680 179.710 ;
        RECT 80.595 179.550 80.885 179.570 ;
        RECT 82.360 179.510 82.680 179.570 ;
        RECT 85.670 179.570 86.345 179.710 ;
        RECT 75.000 179.170 75.320 179.430 ;
        RECT 85.670 179.090 85.810 179.570 ;
        RECT 86.055 179.525 86.345 179.570 ;
        RECT 98.550 179.370 98.690 179.865 ;
        RECT 99.840 179.850 100.160 179.910 ;
        RECT 99.395 179.710 99.685 179.755 ;
        RECT 100.300 179.710 100.620 179.770 ;
        RECT 105.450 179.755 105.590 179.910 ;
        RECT 102.155 179.710 102.445 179.755 ;
        RECT 99.395 179.570 102.445 179.710 ;
        RECT 99.395 179.525 99.685 179.570 ;
        RECT 100.300 179.510 100.620 179.570 ;
        RECT 102.155 179.525 102.445 179.570 ;
        RECT 103.075 179.525 103.365 179.755 ;
        RECT 103.535 179.525 103.825 179.755 ;
        RECT 105.375 179.525 105.665 179.755 ;
        RECT 103.150 179.370 103.290 179.525 ;
        RECT 98.550 179.230 103.290 179.370 ;
        RECT 103.610 179.370 103.750 179.525 ;
        RECT 105.820 179.510 106.140 179.770 ;
        RECT 106.740 179.755 107.060 179.770 ;
        RECT 106.710 179.710 107.060 179.755 ;
        RECT 106.545 179.570 107.060 179.710 ;
        RECT 106.710 179.525 107.060 179.570 ;
        RECT 106.740 179.510 107.060 179.525 ;
        RECT 105.910 179.370 106.050 179.510 ;
        RECT 103.610 179.230 106.050 179.370 ;
        RECT 106.255 179.370 106.545 179.415 ;
        RECT 107.445 179.370 107.735 179.415 ;
        RECT 109.965 179.370 110.255 179.415 ;
        RECT 106.255 179.230 110.255 179.370 ;
        RECT 106.255 179.185 106.545 179.230 ;
        RECT 107.445 179.185 107.735 179.230 ;
        RECT 109.965 179.185 110.255 179.230 ;
        RECT 74.505 179.030 74.795 179.075 ;
        RECT 76.395 179.030 76.685 179.075 ;
        RECT 79.515 179.030 79.805 179.075 ;
        RECT 74.505 178.890 79.805 179.030 ;
        RECT 74.505 178.845 74.795 178.890 ;
        RECT 76.395 178.845 76.685 178.890 ;
        RECT 79.515 178.845 79.805 178.890 ;
        RECT 82.375 179.030 82.665 179.075 ;
        RECT 85.580 179.030 85.900 179.090 ;
        RECT 82.375 178.890 85.900 179.030 ;
        RECT 82.375 178.845 82.665 178.890 ;
        RECT 85.580 178.830 85.900 178.890 ;
        RECT 105.860 179.030 106.150 179.075 ;
        RECT 107.960 179.030 108.250 179.075 ;
        RECT 109.530 179.030 109.820 179.075 ;
        RECT 105.860 178.890 109.820 179.030 ;
        RECT 105.860 178.845 106.150 178.890 ;
        RECT 107.960 178.845 108.250 178.890 ;
        RECT 109.530 178.845 109.820 178.890 ;
        RECT 85.120 178.490 85.440 178.750 ;
        RECT 97.080 178.690 97.400 178.750 ;
        RECT 97.555 178.690 97.845 178.735 ;
        RECT 97.080 178.550 97.845 178.690 ;
        RECT 97.080 178.490 97.400 178.550 ;
        RECT 97.555 178.505 97.845 178.550 ;
        RECT 112.260 178.490 112.580 178.750 ;
        RECT 68.930 177.870 119.550 178.350 ;
        RECT 68.930 172.910 69.410 177.870 ;
        RECT 73.635 177.670 73.925 177.715 ;
        RECT 75.000 177.670 75.320 177.730 ;
        RECT 73.635 177.530 75.320 177.670 ;
        RECT 73.635 177.485 73.925 177.530 ;
        RECT 75.000 177.470 75.320 177.530 ;
        RECT 99.395 177.670 99.685 177.715 ;
        RECT 99.840 177.670 100.160 177.730 ;
        RECT 99.395 177.530 100.160 177.670 ;
        RECT 99.395 177.485 99.685 177.530 ;
        RECT 99.840 177.470 100.160 177.530 ;
        RECT 101.235 177.670 101.525 177.715 ;
        RECT 103.060 177.670 103.380 177.730 ;
        RECT 101.235 177.530 103.380 177.670 ;
        RECT 101.235 177.485 101.525 177.530 ;
        RECT 96.160 177.330 96.480 177.390 ;
        RECT 101.310 177.330 101.450 177.485 ;
        RECT 103.060 177.470 103.380 177.530 ;
        RECT 115.020 177.470 115.340 177.730 ;
        RECT 96.160 177.190 101.450 177.330 ;
        RECT 96.160 177.130 96.480 177.190 ;
        RECT 75.015 176.805 75.305 177.035 ;
        RECT 80.995 176.990 81.285 177.035 ;
        RECT 81.440 176.990 81.760 177.050 ;
        RECT 83.295 176.990 83.585 177.035 ;
        RECT 85.120 176.990 85.440 177.050 ;
        RECT 111.340 176.990 111.660 177.050 ;
        RECT 113.195 176.990 113.485 177.035 ;
        RECT 118.700 176.990 119.020 177.050 ;
        RECT 80.995 176.850 81.760 176.990 ;
        RECT 80.995 176.805 81.285 176.850 ;
        RECT 75.090 176.310 75.230 176.805 ;
        RECT 81.440 176.790 81.760 176.850 ;
        RECT 82.450 176.850 85.440 176.990 ;
        RECT 75.475 176.650 75.765 176.695 ;
        RECT 82.450 176.650 82.590 176.850 ;
        RECT 83.295 176.805 83.585 176.850 ;
        RECT 85.120 176.790 85.440 176.850 ;
        RECT 97.170 176.850 113.485 176.990 ;
        RECT 97.170 176.710 97.310 176.850 ;
        RECT 111.340 176.790 111.660 176.850 ;
        RECT 113.195 176.805 113.485 176.850 ;
        RECT 115.570 176.850 119.020 176.990 ;
        RECT 75.475 176.510 82.590 176.650 ;
        RECT 75.475 176.465 75.765 176.510 ;
        RECT 82.820 176.450 83.140 176.710 ;
        RECT 97.080 176.450 97.400 176.710 ;
        RECT 103.520 176.650 103.840 176.710 ;
        RECT 103.995 176.650 104.285 176.695 ;
        RECT 103.520 176.510 104.285 176.650 ;
        RECT 103.520 176.450 103.840 176.510 ;
        RECT 103.995 176.465 104.285 176.510 ;
        RECT 108.580 176.450 108.900 176.710 ;
        RECT 112.260 176.450 112.580 176.710 ;
        RECT 115.570 176.695 115.710 176.850 ;
        RECT 118.700 176.790 119.020 176.850 ;
        RECT 114.575 176.650 114.865 176.695 ;
        RECT 114.575 176.510 115.250 176.650 ;
        RECT 114.575 176.465 114.865 176.510 ;
        RECT 83.740 176.310 84.060 176.370 ;
        RECT 75.090 176.170 84.060 176.310 ;
        RECT 83.740 176.110 84.060 176.170 ;
        RECT 92.035 176.310 92.325 176.355 ;
        RECT 96.620 176.310 96.940 176.370 ;
        RECT 92.035 176.170 96.940 176.310 ;
        RECT 92.035 176.125 92.325 176.170 ;
        RECT 96.620 176.110 96.940 176.170 ;
        RECT 115.110 176.030 115.250 176.510 ;
        RECT 115.495 176.465 115.785 176.695 ;
        RECT 115.955 176.465 116.245 176.695 ;
        RECT 116.875 176.650 117.165 176.695 ;
        RECT 116.875 176.510 119.850 176.650 ;
        RECT 116.875 176.465 117.165 176.510 ;
        RECT 116.030 176.310 116.170 176.465 ;
        RECT 116.030 176.170 118.010 176.310 ;
        RECT 117.870 176.030 118.010 176.170 ;
        RECT 105.375 175.970 105.665 176.015 ;
        RECT 105.820 175.970 106.140 176.030 ;
        RECT 105.375 175.830 106.140 175.970 ;
        RECT 105.375 175.785 105.665 175.830 ;
        RECT 105.820 175.770 106.140 175.830 ;
        RECT 107.200 175.970 107.520 176.030 ;
        RECT 110.435 175.970 110.725 176.015 ;
        RECT 107.200 175.830 110.725 175.970 ;
        RECT 107.200 175.770 107.520 175.830 ;
        RECT 110.435 175.785 110.725 175.830 ;
        RECT 112.735 175.970 113.025 176.015 ;
        RECT 114.560 175.970 114.880 176.030 ;
        RECT 112.735 175.830 114.880 175.970 ;
        RECT 112.735 175.785 113.025 175.830 ;
        RECT 114.560 175.770 114.880 175.830 ;
        RECT 115.020 175.770 115.340 176.030 ;
        RECT 115.480 175.970 115.800 176.030 ;
        RECT 115.955 175.970 116.245 176.015 ;
        RECT 115.480 175.830 116.245 175.970 ;
        RECT 115.480 175.770 115.800 175.830 ;
        RECT 115.955 175.785 116.245 175.830 ;
        RECT 117.780 175.770 118.100 176.030 ;
        RECT 119.710 175.630 119.850 176.510 ;
        RECT 121.455 175.630 121.935 180.590 ;
        RECT 71.250 175.150 121.935 175.630 ;
        RECT 79.140 174.950 79.460 175.010 ;
        RECT 74.170 174.810 97.770 174.950 ;
        RECT 73.620 174.270 73.940 174.330 ;
        RECT 74.170 174.315 74.310 174.810 ;
        RECT 79.140 174.750 79.460 174.810 ;
        RECT 77.755 174.610 78.405 174.655 ;
        RECT 81.355 174.610 81.645 174.655 ;
        RECT 77.755 174.470 81.645 174.610 ;
        RECT 77.755 174.425 78.405 174.470 ;
        RECT 81.055 174.425 81.645 174.470 ;
        RECT 74.095 174.270 74.385 174.315 ;
        RECT 73.620 174.130 74.385 174.270 ;
        RECT 73.620 174.070 73.940 174.130 ;
        RECT 74.095 174.085 74.385 174.130 ;
        RECT 74.560 174.270 74.850 174.315 ;
        RECT 76.395 174.270 76.685 174.315 ;
        RECT 79.975 174.270 80.265 174.315 ;
        RECT 74.560 174.130 80.265 174.270 ;
        RECT 74.560 174.085 74.850 174.130 ;
        RECT 76.395 174.085 76.685 174.130 ;
        RECT 79.975 174.085 80.265 174.130 ;
        RECT 81.055 174.270 81.345 174.425 ;
        RECT 82.360 174.270 82.680 174.330 ;
        RECT 84.750 174.315 84.890 174.810 ;
        RECT 88.335 174.610 88.985 174.655 ;
        RECT 91.935 174.610 92.225 174.655 ;
        RECT 88.335 174.470 92.225 174.610 ;
        RECT 88.335 174.425 88.985 174.470 ;
        RECT 91.635 174.425 92.225 174.470 ;
        RECT 97.630 174.610 97.770 174.810 ;
        RECT 99.840 174.750 100.160 175.010 ;
        RECT 103.520 174.950 103.840 175.010 ;
        RECT 104.455 174.950 104.745 174.995 ;
        RECT 103.520 174.810 104.745 174.950 ;
        RECT 103.520 174.750 103.840 174.810 ;
        RECT 104.455 174.765 104.745 174.810 ;
        RECT 107.200 174.750 107.520 175.010 ;
        RECT 108.580 174.950 108.900 175.010 ;
        RECT 109.055 174.950 109.345 174.995 ;
        RECT 108.580 174.810 109.345 174.950 ;
        RECT 108.580 174.750 108.900 174.810 ;
        RECT 109.055 174.765 109.345 174.810 ;
        RECT 111.800 174.950 112.120 175.010 ;
        RECT 113.195 174.950 113.485 174.995 ;
        RECT 111.800 174.810 113.485 174.950 ;
        RECT 111.800 174.750 112.120 174.810 ;
        RECT 113.195 174.765 113.485 174.810 ;
        RECT 99.930 174.610 100.070 174.750 ;
        RECT 97.630 174.470 100.070 174.610 ;
        RECT 106.280 174.610 106.600 174.670 ;
        RECT 112.735 174.610 113.025 174.655 ;
        RECT 116.415 174.610 116.705 174.655 ;
        RECT 106.280 174.470 109.730 174.610 ;
        RECT 81.055 174.130 82.680 174.270 ;
        RECT 81.055 174.110 81.345 174.130 ;
        RECT 75.460 173.730 75.780 173.990 ;
        RECT 74.965 173.590 75.255 173.635 ;
        RECT 76.855 173.590 77.145 173.635 ;
        RECT 79.975 173.590 80.265 173.635 ;
        RECT 74.965 173.450 80.265 173.590 ;
        RECT 81.070 173.590 81.210 174.110 ;
        RECT 82.360 174.070 82.680 174.130 ;
        RECT 84.675 174.085 84.965 174.315 ;
        RECT 85.140 174.270 85.430 174.315 ;
        RECT 86.975 174.270 87.265 174.315 ;
        RECT 90.555 174.270 90.845 174.315 ;
        RECT 85.140 174.130 90.845 174.270 ;
        RECT 85.140 174.085 85.430 174.130 ;
        RECT 86.975 174.085 87.265 174.130 ;
        RECT 90.555 174.085 90.845 174.130 ;
        RECT 91.635 174.270 91.925 174.425 ;
        RECT 93.860 174.270 94.180 174.330 ;
        RECT 91.635 174.130 94.180 174.270 ;
        RECT 91.635 174.110 91.925 174.130 ;
        RECT 81.440 173.930 81.760 173.990 ;
        RECT 86.055 173.930 86.345 173.975 ;
        RECT 81.440 173.790 86.345 173.930 ;
        RECT 81.440 173.730 81.760 173.790 ;
        RECT 86.055 173.745 86.345 173.790 ;
        RECT 85.545 173.590 85.835 173.635 ;
        RECT 87.435 173.590 87.725 173.635 ;
        RECT 90.555 173.590 90.845 173.635 ;
        RECT 81.070 173.450 83.510 173.590 ;
        RECT 74.965 173.405 75.255 173.450 ;
        RECT 76.855 173.405 77.145 173.450 ;
        RECT 79.975 173.405 80.265 173.450 ;
        RECT 82.820 173.050 83.140 173.310 ;
        RECT 83.370 173.250 83.510 173.450 ;
        RECT 85.545 173.450 90.845 173.590 ;
        RECT 85.545 173.405 85.835 173.450 ;
        RECT 87.435 173.405 87.725 173.450 ;
        RECT 90.555 173.405 90.845 173.450 ;
        RECT 91.650 173.250 91.790 174.110 ;
        RECT 93.860 174.070 94.180 174.130 ;
        RECT 95.255 174.270 95.545 174.315 ;
        RECT 97.080 174.270 97.400 174.330 ;
        RECT 97.630 174.315 97.770 174.470 ;
        RECT 106.280 174.410 106.600 174.470 ;
        RECT 95.255 174.130 97.400 174.270 ;
        RECT 95.255 174.085 95.545 174.130 ;
        RECT 97.080 174.070 97.400 174.130 ;
        RECT 97.555 174.085 97.845 174.315 ;
        RECT 98.835 174.270 99.125 174.315 ;
        RECT 107.660 174.270 107.980 174.330 ;
        RECT 109.590 174.315 109.730 174.470 ;
        RECT 112.735 174.470 118.010 174.610 ;
        RECT 112.735 174.425 113.025 174.470 ;
        RECT 116.415 174.425 116.705 174.470 ;
        RECT 117.870 174.330 118.010 174.470 ;
        RECT 98.090 174.130 99.125 174.270 ;
        RECT 96.160 173.930 96.480 173.990 ;
        RECT 96.635 173.930 96.925 173.975 ;
        RECT 98.090 173.930 98.230 174.130 ;
        RECT 98.835 174.085 99.125 174.130 ;
        RECT 106.370 174.130 107.980 174.270 ;
        RECT 106.370 173.975 106.510 174.130 ;
        RECT 107.660 174.070 107.980 174.130 ;
        RECT 109.515 174.085 109.805 174.315 ;
        RECT 110.435 174.270 110.725 174.315 ;
        RECT 110.435 174.130 115.250 174.270 ;
        RECT 110.435 174.085 110.725 174.130 ;
        RECT 115.110 173.990 115.250 174.130 ;
        RECT 117.320 174.070 117.640 174.330 ;
        RECT 117.780 174.070 118.100 174.330 ;
        RECT 96.160 173.790 96.925 173.930 ;
        RECT 96.160 173.730 96.480 173.790 ;
        RECT 96.635 173.745 96.925 173.790 ;
        RECT 97.630 173.790 98.230 173.930 ;
        RECT 98.435 173.930 98.725 173.975 ;
        RECT 99.625 173.930 99.915 173.975 ;
        RECT 102.145 173.930 102.435 173.975 ;
        RECT 98.435 173.790 102.435 173.930 ;
        RECT 94.335 173.590 94.625 173.635 ;
        RECT 97.630 173.590 97.770 173.790 ;
        RECT 98.435 173.745 98.725 173.790 ;
        RECT 99.625 173.745 99.915 173.790 ;
        RECT 102.145 173.745 102.435 173.790 ;
        RECT 106.295 173.745 106.585 173.975 ;
        RECT 106.755 173.930 107.045 173.975 ;
        RECT 108.580 173.930 108.900 173.990 ;
        RECT 106.755 173.790 108.900 173.930 ;
        RECT 106.755 173.745 107.045 173.790 ;
        RECT 108.580 173.730 108.900 173.790 ;
        RECT 111.340 173.930 111.660 173.990 ;
        RECT 111.815 173.930 112.105 173.975 ;
        RECT 111.340 173.790 112.105 173.930 ;
        RECT 111.340 173.730 111.660 173.790 ;
        RECT 111.815 173.745 112.105 173.790 ;
        RECT 115.020 173.930 115.340 173.990 ;
        RECT 117.410 173.930 117.550 174.070 ;
        RECT 119.710 173.930 119.850 175.150 ;
        RECT 115.020 173.790 115.710 173.930 ;
        RECT 117.410 173.790 119.850 173.930 ;
        RECT 115.020 173.730 115.340 173.790 ;
        RECT 94.335 173.450 97.770 173.590 ;
        RECT 98.040 173.590 98.330 173.635 ;
        RECT 100.140 173.590 100.430 173.635 ;
        RECT 101.710 173.590 102.000 173.635 ;
        RECT 98.040 173.450 102.000 173.590 ;
        RECT 94.335 173.405 94.625 173.450 ;
        RECT 98.040 173.405 98.330 173.450 ;
        RECT 100.140 173.405 100.430 173.450 ;
        RECT 101.710 173.405 102.000 173.450 ;
        RECT 83.370 173.110 91.790 173.250 ;
        RECT 93.400 173.050 93.720 173.310 ;
        RECT 96.175 173.250 96.465 173.295 ;
        RECT 110.435 173.250 110.725 173.295 ;
        RECT 96.175 173.110 110.725 173.250 ;
        RECT 96.175 173.065 96.465 173.110 ;
        RECT 110.435 173.065 110.725 173.110 ;
        RECT 115.020 173.050 115.340 173.310 ;
        RECT 115.570 173.295 115.710 173.790 ;
        RECT 115.495 173.250 115.785 173.295 ;
        RECT 118.240 173.250 118.560 173.310 ;
        RECT 115.495 173.110 118.560 173.250 ;
        RECT 115.495 173.065 115.785 173.110 ;
        RECT 118.240 173.050 118.560 173.110 ;
        RECT 68.930 172.430 119.550 172.910 ;
        RECT 68.930 167.470 69.410 172.430 ;
        RECT 75.460 172.030 75.780 172.290 ;
        RECT 83.740 172.230 84.060 172.290 ;
        RECT 85.595 172.230 85.885 172.275 ;
        RECT 83.740 172.090 85.885 172.230 ;
        RECT 83.740 172.030 84.060 172.090 ;
        RECT 85.595 172.045 85.885 172.090 ;
        RECT 108.580 172.230 108.900 172.290 ;
        RECT 110.435 172.230 110.725 172.275 ;
        RECT 108.580 172.090 110.725 172.230 ;
        RECT 108.580 172.030 108.900 172.090 ;
        RECT 110.435 172.045 110.725 172.090 ;
        RECT 103.100 171.890 103.390 171.935 ;
        RECT 105.200 171.890 105.490 171.935 ;
        RECT 106.770 171.890 107.060 171.935 ;
        RECT 103.100 171.750 107.060 171.890 ;
        RECT 103.100 171.705 103.390 171.750 ;
        RECT 105.200 171.705 105.490 171.750 ;
        RECT 106.770 171.705 107.060 171.750 ;
        RECT 109.515 171.890 109.805 171.935 ;
        RECT 117.320 171.890 117.640 171.950 ;
        RECT 109.515 171.750 117.640 171.890 ;
        RECT 109.515 171.705 109.805 171.750 ;
        RECT 75.000 171.550 75.320 171.610 ;
        RECT 76.395 171.550 76.685 171.595 ;
        RECT 81.440 171.550 81.760 171.610 ;
        RECT 75.000 171.410 76.685 171.550 ;
        RECT 75.000 171.350 75.320 171.410 ;
        RECT 76.395 171.365 76.685 171.410 ;
        RECT 79.460 171.410 81.760 171.550 ;
        RECT 76.855 171.210 77.145 171.255 ;
        RECT 79.460 171.210 79.600 171.410 ;
        RECT 81.440 171.350 81.760 171.410 ;
        RECT 82.360 171.550 82.680 171.610 ;
        RECT 90.655 171.550 90.945 171.595 ;
        RECT 82.360 171.410 90.945 171.550 ;
        RECT 82.360 171.350 82.680 171.410 ;
        RECT 90.655 171.365 90.945 171.410 ;
        RECT 92.035 171.550 92.325 171.595 ;
        RECT 93.400 171.550 93.720 171.610 ;
        RECT 113.270 171.595 113.410 171.750 ;
        RECT 117.320 171.690 117.640 171.750 ;
        RECT 92.035 171.410 93.720 171.550 ;
        RECT 92.035 171.365 92.325 171.410 ;
        RECT 93.400 171.350 93.720 171.410 ;
        RECT 103.495 171.550 103.785 171.595 ;
        RECT 104.685 171.550 104.975 171.595 ;
        RECT 107.205 171.550 107.495 171.595 ;
        RECT 103.495 171.410 107.495 171.550 ;
        RECT 103.495 171.365 103.785 171.410 ;
        RECT 104.685 171.365 104.975 171.410 ;
        RECT 107.205 171.365 107.495 171.410 ;
        RECT 113.195 171.365 113.485 171.595 ;
        RECT 115.020 171.550 115.340 171.610 ;
        RECT 116.875 171.550 117.165 171.595 ;
        RECT 115.020 171.410 117.165 171.550 ;
        RECT 115.020 171.350 115.340 171.410 ;
        RECT 116.875 171.365 117.165 171.410 ;
        RECT 82.820 171.210 83.140 171.270 ;
        RECT 84.675 171.210 84.965 171.255 ;
        RECT 76.855 171.070 79.600 171.210 ;
        RECT 81.530 171.070 84.965 171.210 ;
        RECT 76.855 171.025 77.145 171.070 ;
        RECT 81.530 170.590 81.670 171.070 ;
        RECT 82.820 171.010 83.140 171.070 ;
        RECT 84.675 171.025 84.965 171.070 ;
        RECT 102.615 171.210 102.905 171.255 ;
        RECT 102.615 171.070 108.350 171.210 ;
        RECT 102.615 171.025 102.905 171.070 ;
        RECT 86.500 170.870 86.820 170.930 ;
        RECT 92.495 170.870 92.785 170.915 ;
        RECT 86.500 170.730 92.785 170.870 ;
        RECT 86.500 170.670 86.820 170.730 ;
        RECT 92.495 170.685 92.785 170.730 ;
        RECT 103.060 170.870 103.380 170.930 ;
        RECT 103.840 170.870 104.130 170.915 ;
        RECT 103.060 170.730 104.130 170.870 ;
        RECT 103.060 170.670 103.380 170.730 ;
        RECT 103.840 170.685 104.130 170.730 ;
        RECT 108.210 170.590 108.350 171.070 ;
        RECT 81.440 170.330 81.760 170.590 ;
        RECT 96.620 170.530 96.940 170.590 ;
        RECT 98.935 170.530 99.225 170.575 ;
        RECT 96.620 170.390 99.225 170.530 ;
        RECT 96.620 170.330 96.940 170.390 ;
        RECT 98.935 170.345 99.225 170.390 ;
        RECT 108.120 170.330 108.440 170.590 ;
        RECT 114.100 170.330 114.420 170.590 ;
        RECT 121.455 170.190 121.935 175.150 ;
        RECT 71.250 169.710 121.935 170.190 ;
        RECT 103.060 169.510 103.380 169.570 ;
        RECT 104.455 169.510 104.745 169.555 ;
        RECT 103.060 169.370 104.745 169.510 ;
        RECT 103.060 169.310 103.380 169.370 ;
        RECT 104.455 169.325 104.745 169.370 ;
        RECT 105.820 169.310 106.140 169.570 ;
        RECT 110.435 169.325 110.725 169.555 ;
        RECT 85.580 168.630 85.900 168.890 ;
        RECT 88.815 168.830 89.105 168.875 ;
        RECT 90.180 168.830 90.500 168.890 ;
        RECT 88.815 168.690 90.500 168.830 ;
        RECT 88.815 168.645 89.105 168.690 ;
        RECT 90.180 168.630 90.500 168.690 ;
        RECT 93.860 168.830 94.180 168.890 ;
        RECT 97.555 168.830 97.845 168.875 ;
        RECT 93.860 168.690 97.845 168.830 ;
        RECT 93.860 168.630 94.180 168.690 ;
        RECT 97.555 168.645 97.845 168.690 ;
        RECT 105.375 168.830 105.665 168.875 ;
        RECT 105.910 168.830 106.050 169.310 ;
        RECT 110.510 169.170 110.650 169.325 ;
        RECT 114.100 169.310 114.420 169.570 ;
        RECT 117.780 169.310 118.100 169.570 ;
        RECT 112.120 169.170 112.410 169.215 ;
        RECT 110.510 169.030 112.410 169.170 ;
        RECT 112.120 168.985 112.410 169.030 ;
        RECT 105.375 168.690 106.050 168.830 ;
        RECT 107.660 168.830 107.980 168.890 ;
        RECT 108.595 168.830 108.885 168.875 ;
        RECT 114.190 168.830 114.330 169.310 ;
        RECT 107.660 168.690 108.885 168.830 ;
        RECT 105.375 168.645 105.665 168.690 ;
        RECT 107.660 168.630 107.980 168.690 ;
        RECT 108.595 168.645 108.885 168.690 ;
        RECT 109.130 168.690 114.330 168.830 ;
        RECT 82.360 168.290 82.680 168.550 ;
        RECT 83.740 168.490 84.060 168.550 ;
        RECT 109.130 168.535 109.270 168.690 ;
        RECT 85.135 168.490 85.425 168.535 ;
        RECT 88.355 168.490 88.645 168.535 ;
        RECT 83.740 168.350 85.425 168.490 ;
        RECT 83.740 168.290 84.060 168.350 ;
        RECT 85.135 168.305 85.425 168.350 ;
        RECT 86.590 168.350 88.645 168.490 ;
        RECT 82.450 168.150 82.590 168.290 ;
        RECT 86.590 168.150 86.730 168.350 ;
        RECT 88.355 168.305 88.645 168.350 ;
        RECT 91.115 168.305 91.405 168.535 ;
        RECT 109.055 168.305 109.345 168.535 ;
        RECT 110.895 168.305 111.185 168.535 ;
        RECT 111.775 168.490 112.065 168.535 ;
        RECT 112.965 168.490 113.255 168.535 ;
        RECT 115.485 168.490 115.775 168.535 ;
        RECT 111.775 168.350 115.775 168.490 ;
        RECT 111.775 168.305 112.065 168.350 ;
        RECT 112.965 168.305 113.255 168.350 ;
        RECT 115.485 168.305 115.775 168.350 ;
        RECT 82.450 168.010 86.730 168.150 ;
        RECT 87.435 168.150 87.725 168.195 ;
        RECT 91.190 168.150 91.330 168.305 ;
        RECT 110.970 168.150 111.110 168.305 ;
        RECT 87.435 168.010 91.330 168.150 ;
        RECT 108.210 168.010 111.110 168.150 ;
        RECT 111.380 168.150 111.670 168.195 ;
        RECT 113.480 168.150 113.770 168.195 ;
        RECT 115.050 168.150 115.340 168.195 ;
        RECT 111.380 168.010 115.340 168.150 ;
        RECT 87.435 167.965 87.725 168.010 ;
        RECT 108.210 167.870 108.350 168.010 ;
        RECT 111.380 167.965 111.670 168.010 ;
        RECT 113.480 167.965 113.770 168.010 ;
        RECT 115.050 167.965 115.340 168.010 ;
        RECT 90.655 167.810 90.945 167.855 ;
        RECT 93.860 167.810 94.180 167.870 ;
        RECT 90.655 167.670 94.180 167.810 ;
        RECT 90.655 167.625 90.945 167.670 ;
        RECT 93.860 167.610 94.180 167.670 ;
        RECT 94.335 167.810 94.625 167.855 ;
        RECT 94.780 167.810 95.100 167.870 ;
        RECT 94.335 167.670 95.100 167.810 ;
        RECT 94.335 167.625 94.625 167.670 ;
        RECT 94.780 167.610 95.100 167.670 ;
        RECT 95.700 167.810 96.020 167.870 ;
        RECT 98.475 167.810 98.765 167.855 ;
        RECT 95.700 167.670 98.765 167.810 ;
        RECT 95.700 167.610 96.020 167.670 ;
        RECT 98.475 167.625 98.765 167.670 ;
        RECT 108.120 167.610 108.440 167.870 ;
        RECT 68.930 166.990 119.550 167.470 ;
        RECT 68.930 162.030 69.410 166.990 ;
        RECT 75.000 166.590 75.320 166.850 ;
        RECT 102.155 166.790 102.445 166.835 ;
        RECT 106.280 166.790 106.600 166.850 ;
        RECT 107.675 166.790 107.965 166.835 ;
        RECT 102.155 166.650 107.965 166.790 ;
        RECT 102.155 166.605 102.445 166.650 ;
        RECT 106.280 166.590 106.600 166.650 ;
        RECT 107.675 166.605 107.965 166.650 ;
        RECT 115.480 166.590 115.800 166.850 ;
        RECT 77.775 166.265 78.065 166.495 ;
        RECT 94.285 166.450 94.575 166.495 ;
        RECT 96.175 166.450 96.465 166.495 ;
        RECT 99.295 166.450 99.585 166.495 ;
        RECT 94.285 166.310 99.585 166.450 ;
        RECT 94.285 166.265 94.575 166.310 ;
        RECT 96.175 166.265 96.465 166.310 ;
        RECT 99.295 166.265 99.585 166.310 ;
        RECT 76.855 166.110 77.145 166.155 ;
        RECT 77.850 166.110 77.990 166.265 ;
        RECT 76.855 165.970 77.990 166.110 ;
        RECT 80.075 166.110 80.365 166.155 ;
        RECT 81.440 166.110 81.760 166.170 ;
        RECT 80.075 165.970 81.760 166.110 ;
        RECT 76.855 165.925 77.145 165.970 ;
        RECT 80.075 165.925 80.365 165.970 ;
        RECT 81.440 165.910 81.760 165.970 ;
        RECT 82.360 165.910 82.680 166.170 ;
        RECT 83.755 166.110 84.045 166.155 ;
        RECT 86.055 166.110 86.345 166.155 ;
        RECT 83.755 165.970 86.345 166.110 ;
        RECT 83.755 165.925 84.045 165.970 ;
        RECT 86.055 165.925 86.345 165.970 ;
        RECT 94.780 165.910 95.100 166.170 ;
        RECT 115.570 166.110 115.710 166.590 ;
        RECT 115.570 165.970 116.630 166.110 ;
        RECT 76.395 165.770 76.685 165.815 ;
        RECT 79.615 165.770 79.905 165.815 ;
        RECT 80.980 165.770 81.300 165.830 ;
        RECT 76.395 165.630 77.070 165.770 ;
        RECT 76.395 165.585 76.685 165.630 ;
        RECT 76.930 165.150 77.070 165.630 ;
        RECT 79.615 165.630 81.300 165.770 ;
        RECT 79.615 165.585 79.905 165.630 ;
        RECT 80.980 165.570 81.300 165.630 ;
        RECT 81.915 165.770 82.205 165.815 ;
        RECT 85.580 165.770 85.900 165.830 ;
        RECT 92.955 165.770 93.245 165.815 ;
        RECT 81.915 165.630 93.245 165.770 ;
        RECT 81.915 165.585 82.205 165.630 ;
        RECT 85.580 165.570 85.900 165.630 ;
        RECT 92.955 165.585 93.245 165.630 ;
        RECT 93.415 165.585 93.705 165.815 ;
        RECT 93.880 165.770 94.170 165.815 ;
        RECT 95.715 165.770 96.005 165.815 ;
        RECT 99.295 165.770 99.585 165.815 ;
        RECT 93.880 165.630 99.585 165.770 ;
        RECT 93.880 165.585 94.170 165.630 ;
        RECT 95.715 165.585 96.005 165.630 ;
        RECT 99.295 165.585 99.585 165.630 ;
        RECT 93.490 165.430 93.630 165.585 ;
        RECT 100.375 165.475 100.665 165.790 ;
        RECT 109.055 165.770 109.345 165.815 ;
        RECT 109.055 165.630 110.650 165.770 ;
        RECT 109.055 165.585 109.345 165.630 ;
        RECT 97.075 165.430 97.725 165.475 ;
        RECT 100.375 165.430 100.965 165.475 ;
        RECT 93.490 165.290 94.090 165.430 ;
        RECT 93.950 165.150 94.090 165.290 ;
        RECT 95.790 165.290 100.965 165.430 ;
        RECT 95.790 165.150 95.930 165.290 ;
        RECT 97.075 165.245 97.725 165.290 ;
        RECT 100.675 165.245 100.965 165.290 ;
        RECT 110.510 165.150 110.650 165.630 ;
        RECT 114.560 165.570 114.880 165.830 ;
        RECT 116.490 165.815 116.630 165.970 ;
        RECT 115.495 165.585 115.785 165.815 ;
        RECT 116.415 165.585 116.705 165.815 ;
        RECT 115.570 165.430 115.710 165.585 ;
        RECT 118.240 165.430 118.560 165.490 ;
        RECT 115.570 165.290 118.560 165.430 ;
        RECT 118.240 165.230 118.560 165.290 ;
        RECT 76.840 164.890 77.160 165.150 ;
        RECT 89.260 164.890 89.580 165.150 ;
        RECT 90.180 165.090 90.500 165.150 ;
        RECT 92.035 165.090 92.325 165.135 ;
        RECT 90.180 164.950 92.325 165.090 ;
        RECT 90.180 164.890 90.500 164.950 ;
        RECT 92.035 164.905 92.325 164.950 ;
        RECT 93.860 164.890 94.180 165.150 ;
        RECT 95.700 164.890 96.020 165.150 ;
        RECT 106.740 164.890 107.060 165.150 ;
        RECT 110.420 164.890 110.740 165.150 ;
        RECT 111.800 164.890 112.120 165.150 ;
        RECT 115.020 165.090 115.340 165.150 ;
        RECT 115.495 165.090 115.785 165.135 ;
        RECT 115.020 164.950 115.785 165.090 ;
        RECT 115.020 164.890 115.340 164.950 ;
        RECT 115.495 164.905 115.785 164.950 ;
        RECT 121.455 164.750 121.935 169.710 ;
        RECT 71.250 164.270 121.935 164.750 ;
        RECT 85.580 163.870 85.900 164.130 ;
        RECT 89.260 164.070 89.580 164.130 ;
        RECT 95.700 164.070 96.020 164.130 ;
        RECT 89.260 163.930 93.170 164.070 ;
        RECT 89.260 163.870 89.580 163.930 ;
        RECT 93.030 163.775 93.170 163.930 ;
        RECT 95.700 163.930 99.610 164.070 ;
        RECT 95.700 163.870 96.020 163.930 ;
        RECT 79.135 163.730 79.785 163.775 ;
        RECT 82.735 163.730 83.025 163.775 ;
        RECT 79.135 163.590 83.025 163.730 ;
        RECT 79.135 163.545 79.785 163.590 ;
        RECT 82.435 163.545 83.025 163.590 ;
        RECT 87.075 163.730 87.365 163.775 ;
        RECT 90.315 163.730 90.965 163.775 ;
        RECT 87.075 163.590 90.965 163.730 ;
        RECT 87.075 163.545 87.665 163.590 ;
        RECT 90.315 163.545 90.965 163.590 ;
        RECT 92.955 163.545 93.245 163.775 ;
        RECT 94.320 163.730 94.640 163.790 ;
        RECT 98.935 163.730 99.225 163.775 ;
        RECT 94.320 163.590 99.225 163.730 ;
        RECT 99.470 163.730 99.610 163.930 ;
        RECT 101.215 163.730 101.865 163.775 ;
        RECT 104.815 163.730 105.105 163.775 ;
        RECT 99.470 163.590 105.105 163.730 ;
        RECT 75.940 163.390 76.230 163.435 ;
        RECT 77.775 163.390 78.065 163.435 ;
        RECT 81.355 163.390 81.645 163.435 ;
        RECT 75.940 163.250 81.645 163.390 ;
        RECT 75.940 163.205 76.230 163.250 ;
        RECT 77.775 163.205 78.065 163.250 ;
        RECT 81.355 163.205 81.645 163.250 ;
        RECT 82.435 163.390 82.725 163.545 ;
        RECT 87.375 163.390 87.665 163.545 ;
        RECT 94.320 163.530 94.640 163.590 ;
        RECT 98.935 163.545 99.225 163.590 ;
        RECT 101.215 163.545 101.865 163.590 ;
        RECT 104.515 163.545 105.105 163.590 ;
        RECT 109.470 163.730 109.760 163.775 ;
        RECT 111.800 163.730 112.120 163.790 ;
        RECT 109.470 163.590 112.120 163.730 ;
        RECT 109.470 163.545 109.760 163.590 ;
        RECT 82.435 163.250 87.665 163.390 ;
        RECT 82.435 163.230 82.725 163.250 ;
        RECT 75.460 162.850 75.780 163.110 ;
        RECT 76.840 163.050 77.160 163.110 ;
        RECT 79.140 163.050 79.460 163.110 ;
        RECT 76.840 162.910 79.460 163.050 ;
        RECT 76.840 162.850 77.160 162.910 ;
        RECT 79.140 162.850 79.460 162.910 ;
        RECT 76.345 162.710 76.635 162.755 ;
        RECT 78.235 162.710 78.525 162.755 ;
        RECT 81.355 162.710 81.645 162.755 ;
        RECT 76.345 162.570 81.645 162.710 ;
        RECT 76.345 162.525 76.635 162.570 ;
        RECT 78.235 162.525 78.525 162.570 ;
        RECT 81.355 162.525 81.645 162.570 ;
        RECT 82.910 162.430 83.050 163.250 ;
        RECT 87.375 163.230 87.665 163.250 ;
        RECT 88.455 163.390 88.745 163.435 ;
        RECT 92.035 163.390 92.325 163.435 ;
        RECT 93.870 163.390 94.160 163.435 ;
        RECT 88.455 163.250 94.160 163.390 ;
        RECT 88.455 163.205 88.745 163.250 ;
        RECT 92.035 163.205 92.325 163.250 ;
        RECT 93.870 163.205 94.160 163.250 ;
        RECT 98.020 163.390 98.310 163.435 ;
        RECT 99.855 163.390 100.145 163.435 ;
        RECT 103.435 163.390 103.725 163.435 ;
        RECT 98.020 163.250 103.725 163.390 ;
        RECT 98.020 163.205 98.310 163.250 ;
        RECT 99.855 163.205 100.145 163.250 ;
        RECT 103.435 163.205 103.725 163.250 ;
        RECT 104.515 163.230 104.805 163.545 ;
        RECT 111.800 163.530 112.120 163.590 ;
        RECT 94.335 163.050 94.625 163.095 ;
        RECT 97.555 163.050 97.845 163.095 ;
        RECT 93.950 162.910 97.845 163.050 ;
        RECT 88.455 162.710 88.745 162.755 ;
        RECT 91.575 162.710 91.865 162.755 ;
        RECT 93.465 162.710 93.755 162.755 ;
        RECT 88.455 162.570 93.755 162.710 ;
        RECT 88.455 162.525 88.745 162.570 ;
        RECT 91.575 162.525 91.865 162.570 ;
        RECT 93.465 162.525 93.755 162.570 ;
        RECT 93.950 162.430 94.090 162.910 ;
        RECT 94.335 162.865 94.625 162.910 ;
        RECT 97.555 162.865 97.845 162.910 ;
        RECT 108.120 162.850 108.440 163.110 ;
        RECT 109.015 163.050 109.305 163.095 ;
        RECT 110.205 163.050 110.495 163.095 ;
        RECT 112.725 163.050 113.015 163.095 ;
        RECT 109.015 162.910 113.015 163.050 ;
        RECT 109.015 162.865 109.305 162.910 ;
        RECT 110.205 162.865 110.495 162.910 ;
        RECT 112.725 162.865 113.015 162.910 ;
        RECT 98.425 162.710 98.715 162.755 ;
        RECT 100.315 162.710 100.605 162.755 ;
        RECT 103.435 162.710 103.725 162.755 ;
        RECT 98.425 162.570 103.725 162.710 ;
        RECT 98.425 162.525 98.715 162.570 ;
        RECT 100.315 162.525 100.605 162.570 ;
        RECT 103.435 162.525 103.725 162.570 ;
        RECT 108.620 162.710 108.910 162.755 ;
        RECT 110.720 162.710 111.010 162.755 ;
        RECT 112.290 162.710 112.580 162.755 ;
        RECT 108.620 162.570 112.580 162.710 ;
        RECT 108.620 162.525 108.910 162.570 ;
        RECT 110.720 162.525 111.010 162.570 ;
        RECT 112.290 162.525 112.580 162.570 ;
        RECT 82.820 162.170 83.140 162.430 ;
        RECT 84.200 162.170 84.520 162.430 ;
        RECT 93.860 162.170 94.180 162.430 ;
        RECT 106.295 162.370 106.585 162.415 ;
        RECT 109.500 162.370 109.820 162.430 ;
        RECT 106.295 162.230 109.820 162.370 ;
        RECT 106.295 162.185 106.585 162.230 ;
        RECT 109.500 162.170 109.820 162.230 ;
        RECT 115.020 162.170 115.340 162.430 ;
        RECT 68.930 161.550 119.550 162.030 ;
        RECT 68.930 156.590 69.410 161.550 ;
        RECT 84.200 161.150 84.520 161.410 ;
        RECT 106.280 161.350 106.600 161.410 ;
        RECT 111.815 161.350 112.105 161.395 ;
        RECT 106.280 161.210 112.105 161.350 ;
        RECT 106.280 161.150 106.600 161.210 ;
        RECT 111.815 161.165 112.105 161.210 ;
        RECT 114.115 161.350 114.405 161.395 ;
        RECT 114.560 161.350 114.880 161.410 ;
        RECT 114.115 161.210 114.880 161.350 ;
        RECT 114.115 161.165 114.405 161.210 ;
        RECT 114.560 161.150 114.880 161.210 ;
        RECT 84.290 160.670 84.430 161.150 ;
        RECT 102.600 161.010 102.920 161.070 ;
        RECT 112.275 161.010 112.565 161.055 ;
        RECT 102.600 160.870 112.565 161.010 ;
        RECT 102.600 160.810 102.920 160.870 ;
        RECT 112.275 160.825 112.565 160.870 ;
        RECT 86.515 160.670 86.805 160.715 ;
        RECT 111.355 160.670 111.645 160.715 ;
        RECT 84.290 160.530 86.805 160.670 ;
        RECT 86.515 160.485 86.805 160.530 ;
        RECT 109.590 160.530 111.645 160.670 ;
        RECT 109.590 160.390 109.730 160.530 ;
        RECT 111.355 160.485 111.645 160.530 ;
        RECT 115.020 160.670 115.340 160.730 ;
        RECT 117.335 160.670 117.625 160.715 ;
        RECT 115.020 160.530 117.625 160.670 ;
        RECT 115.020 160.470 115.340 160.530 ;
        RECT 117.335 160.485 117.625 160.530 ;
        RECT 87.895 160.145 88.185 160.375 ;
        RECT 87.970 159.710 88.110 160.145 ;
        RECT 102.140 160.130 102.460 160.390 ;
        RECT 103.060 160.330 103.380 160.390 ;
        RECT 105.835 160.330 106.125 160.375 ;
        RECT 103.060 160.190 106.125 160.330 ;
        RECT 103.060 160.130 103.380 160.190 ;
        RECT 105.835 160.145 106.125 160.190 ;
        RECT 108.580 160.130 108.900 160.390 ;
        RECT 109.500 160.130 109.820 160.390 ;
        RECT 110.420 160.130 110.740 160.390 ;
        RECT 112.735 160.330 113.025 160.375 ;
        RECT 114.575 160.330 114.865 160.375 ;
        RECT 112.735 160.190 114.865 160.330 ;
        RECT 112.735 160.145 113.025 160.190 ;
        RECT 114.575 160.145 114.865 160.190 ;
        RECT 87.880 159.450 88.200 159.710 ;
        RECT 103.520 159.650 103.840 159.710 ;
        RECT 105.375 159.650 105.665 159.695 ;
        RECT 103.520 159.510 105.665 159.650 ;
        RECT 103.520 159.450 103.840 159.510 ;
        RECT 105.375 159.465 105.665 159.510 ;
        RECT 121.455 159.310 121.935 164.270 ;
        RECT 71.250 158.830 121.935 159.310 ;
        RECT 101.695 158.630 101.985 158.675 ;
        RECT 102.140 158.630 102.460 158.690 ;
        RECT 101.695 158.490 102.460 158.630 ;
        RECT 101.695 158.445 101.985 158.490 ;
        RECT 102.140 158.430 102.460 158.490 ;
        RECT 106.295 158.630 106.585 158.675 ;
        RECT 106.295 158.490 115.710 158.630 ;
        RECT 106.295 158.445 106.585 158.490 ;
        RECT 82.820 158.290 83.140 158.350 ;
        RECT 95.700 158.290 96.020 158.350 ;
        RECT 82.820 158.150 96.020 158.290 ;
        RECT 82.820 158.090 83.140 158.150 ;
        RECT 95.700 158.090 96.020 158.150 ;
        RECT 107.670 158.290 107.960 158.335 ;
        RECT 108.590 158.290 108.880 158.335 ;
        RECT 114.110 158.290 114.400 158.335 ;
        RECT 107.670 158.150 114.400 158.290 ;
        RECT 107.670 158.105 107.960 158.150 ;
        RECT 108.590 158.105 108.880 158.150 ;
        RECT 114.110 158.105 114.400 158.150 ;
        RECT 82.360 157.750 82.680 158.010 ;
        RECT 86.515 157.950 86.805 157.995 ;
        RECT 82.910 157.810 86.805 157.950 ;
        RECT 82.910 157.655 83.050 157.810 ;
        RECT 86.515 157.765 86.805 157.810 ;
        RECT 88.815 157.950 89.105 157.995 ;
        RECT 93.400 157.950 93.720 158.010 ;
        RECT 88.815 157.810 93.720 157.950 ;
        RECT 88.815 157.765 89.105 157.810 ;
        RECT 82.835 157.425 83.125 157.655 ;
        RECT 84.215 157.610 84.505 157.655 ;
        RECT 85.580 157.610 85.900 157.670 ;
        RECT 84.215 157.470 85.900 157.610 ;
        RECT 84.215 157.425 84.505 157.470 ;
        RECT 85.580 157.410 85.900 157.470 ;
        RECT 86.055 157.425 86.345 157.655 ;
        RECT 86.590 157.610 86.730 157.765 ;
        RECT 93.400 157.750 93.720 157.810 ;
        RECT 103.060 157.750 103.380 158.010 ;
        RECT 103.535 157.765 103.825 157.995 ;
        RECT 105.375 157.765 105.665 157.995 ;
        RECT 107.165 157.950 107.455 157.995 ;
        RECT 109.005 157.950 109.295 157.995 ;
        RECT 107.165 157.810 109.295 157.950 ;
        RECT 107.165 157.765 107.455 157.810 ;
        RECT 109.005 157.765 109.295 157.810 ;
        RECT 87.880 157.610 88.200 157.670 ;
        RECT 88.355 157.610 88.645 157.655 ;
        RECT 86.590 157.470 88.645 157.610 ;
        RECT 86.130 157.270 86.270 157.425 ;
        RECT 87.880 157.410 88.200 157.470 ;
        RECT 88.355 157.425 88.645 157.470 ;
        RECT 90.655 157.610 90.945 157.655 ;
        RECT 91.575 157.610 91.865 157.655 ;
        RECT 103.610 157.610 103.750 157.765 ;
        RECT 90.655 157.470 91.865 157.610 ;
        RECT 90.655 157.425 90.945 157.470 ;
        RECT 91.575 157.425 91.865 157.470 ;
        RECT 103.150 157.470 103.750 157.610 ;
        RECT 103.995 157.610 104.285 157.655 ;
        RECT 104.900 157.610 105.220 157.670 ;
        RECT 103.995 157.470 105.220 157.610 ;
        RECT 90.180 157.270 90.500 157.330 ;
        RECT 79.460 157.130 84.890 157.270 ;
        RECT 86.130 157.130 90.500 157.270 ;
        RECT 79.460 156.990 79.600 157.130 ;
        RECT 79.140 156.790 79.600 156.990 ;
        RECT 84.750 156.975 84.890 157.130 ;
        RECT 90.180 157.070 90.500 157.130 ;
        RECT 102.600 157.270 102.920 157.330 ;
        RECT 103.150 157.270 103.290 157.470 ;
        RECT 103.995 157.425 104.285 157.470 ;
        RECT 104.900 157.410 105.220 157.470 ;
        RECT 105.450 157.270 105.590 157.765 ;
        RECT 109.500 157.750 109.820 158.010 ;
        RECT 111.350 157.950 111.640 157.995 ;
        RECT 113.190 157.950 113.480 157.995 ;
        RECT 111.350 157.810 113.480 157.950 ;
        RECT 111.350 157.765 111.640 157.810 ;
        RECT 113.190 157.765 113.480 157.810 ;
        RECT 114.575 157.950 114.865 157.995 ;
        RECT 115.020 157.950 115.340 158.010 ;
        RECT 114.575 157.810 115.340 157.950 ;
        RECT 115.570 157.950 115.710 158.490 ;
        RECT 118.700 157.950 119.020 158.010 ;
        RECT 115.570 157.810 119.020 157.950 ;
        RECT 114.575 157.765 114.865 157.810 ;
        RECT 115.020 157.750 115.340 157.810 ;
        RECT 118.700 157.750 119.020 157.810 ;
        RECT 108.580 157.610 108.900 157.670 ;
        RECT 110.205 157.610 110.495 157.655 ;
        RECT 108.580 157.470 110.495 157.610 ;
        RECT 108.580 157.410 108.900 157.470 ;
        RECT 110.205 157.425 110.495 157.470 ;
        RECT 110.880 157.410 111.200 157.670 ;
        RECT 115.480 157.410 115.800 157.670 ;
        RECT 102.600 157.130 103.290 157.270 ;
        RECT 104.070 157.130 105.590 157.270 ;
        RECT 102.600 157.070 102.920 157.130 ;
        RECT 79.140 156.730 79.460 156.790 ;
        RECT 84.675 156.745 84.965 156.975 ;
        RECT 94.320 156.930 94.640 156.990 ;
        RECT 94.795 156.930 95.085 156.975 ;
        RECT 94.320 156.790 95.085 156.930 ;
        RECT 94.320 156.730 94.640 156.790 ;
        RECT 94.795 156.745 95.085 156.790 ;
        RECT 103.060 156.930 103.380 156.990 ;
        RECT 104.070 156.930 104.210 157.130 ;
        RECT 103.060 156.790 104.210 156.930 ;
        RECT 103.060 156.730 103.380 156.790 ;
        RECT 104.440 156.730 104.760 156.990 ;
        RECT 105.450 156.930 105.590 157.130 ;
        RECT 108.085 157.270 108.375 157.315 ;
        RECT 111.315 157.270 111.605 157.315 ;
        RECT 108.085 157.130 111.605 157.270 ;
        RECT 108.085 157.085 108.375 157.130 ;
        RECT 111.315 157.085 111.605 157.130 ;
        RECT 112.275 157.085 112.565 157.315 ;
        RECT 110.420 156.930 110.740 156.990 ;
        RECT 112.350 156.930 112.490 157.085 ;
        RECT 105.450 156.790 112.490 156.930 ;
        RECT 110.420 156.730 110.740 156.790 ;
        RECT 68.930 156.110 119.550 156.590 ;
        RECT 17.610 152.920 17.985 153.265 ;
        RECT 20.630 153.205 20.965 153.285 ;
        RECT 19.810 153.005 20.965 153.205 ;
        RECT 17.695 150.735 17.885 152.920 ;
        RECT 18.930 151.165 19.160 152.165 ;
        RECT 19.370 151.165 19.600 152.165 ;
        RECT 19.810 151.165 20.040 153.005 ;
        RECT 20.630 152.940 20.965 153.005 ;
        RECT 20.440 151.165 20.670 152.165 ;
        RECT 20.880 151.165 21.110 152.165 ;
        RECT 21.320 151.460 21.550 152.165 ;
        RECT 21.320 151.290 22.470 151.460 ;
        RECT 21.320 151.165 21.550 151.290 ;
        RECT 18.960 150.735 19.130 151.165 ;
        RECT 17.695 150.570 19.140 150.735 ;
        RECT 14.840 147.275 16.515 148.550 ;
        RECT 10.665 141.075 17.380 141.245 ;
        RECT 10.665 124.405 10.835 141.075 ;
        RECT 17.210 136.640 17.380 141.075 ;
        RECT 18.960 139.445 19.130 150.570 ;
        RECT 19.840 147.925 20.010 151.165 ;
        RECT 20.470 150.490 20.640 151.165 ;
        RECT 21.100 150.490 21.330 150.550 ;
        RECT 20.470 150.320 21.330 150.490 ;
        RECT 20.470 150.135 20.640 150.320 ;
        RECT 21.100 150.260 21.330 150.320 ;
        RECT 20.425 149.815 20.685 150.135 ;
        RECT 19.600 147.505 20.050 147.925 ;
        RECT 19.840 140.735 20.010 147.505 ;
        RECT 22.300 144.220 22.470 151.290 ;
        RECT 68.930 151.150 69.410 156.110 ;
        RECT 82.360 155.910 82.680 155.970 ;
        RECT 88.355 155.910 88.645 155.955 ;
        RECT 82.360 155.770 88.645 155.910 ;
        RECT 82.360 155.710 82.680 155.770 ;
        RECT 88.355 155.725 88.645 155.770 ;
        RECT 93.350 155.910 93.640 155.955 ;
        RECT 94.320 155.910 94.640 155.970 ;
        RECT 93.350 155.770 94.640 155.910 ;
        RECT 93.350 155.725 93.640 155.770 ;
        RECT 94.320 155.710 94.640 155.770 ;
        RECT 100.775 155.910 101.065 155.955 ;
        RECT 103.060 155.910 103.380 155.970 ;
        RECT 100.775 155.770 103.380 155.910 ;
        RECT 100.775 155.725 101.065 155.770 ;
        RECT 103.060 155.710 103.380 155.770 ;
        RECT 104.440 155.910 104.760 155.970 ;
        RECT 108.135 155.910 108.425 155.955 ;
        RECT 108.580 155.910 108.900 155.970 ;
        RECT 104.440 155.770 106.970 155.910 ;
        RECT 104.440 155.710 104.760 155.770 ;
        RECT 106.830 155.630 106.970 155.770 ;
        RECT 108.135 155.770 108.900 155.910 ;
        RECT 108.135 155.725 108.425 155.770 ;
        RECT 108.580 155.710 108.900 155.770 ;
        RECT 115.480 155.910 115.800 155.970 ;
        RECT 117.780 155.910 118.100 155.970 ;
        RECT 115.480 155.770 118.100 155.910 ;
        RECT 115.480 155.710 115.800 155.770 ;
        RECT 117.780 155.710 118.100 155.770 ;
        RECT 74.505 155.570 74.795 155.615 ;
        RECT 76.395 155.570 76.685 155.615 ;
        RECT 79.515 155.570 79.805 155.615 ;
        RECT 74.505 155.430 79.805 155.570 ;
        RECT 74.505 155.385 74.795 155.430 ;
        RECT 76.395 155.385 76.685 155.430 ;
        RECT 79.515 155.385 79.805 155.430 ;
        RECT 92.905 155.570 93.195 155.615 ;
        RECT 94.795 155.570 95.085 155.615 ;
        RECT 97.915 155.570 98.205 155.615 ;
        RECT 92.905 155.430 98.205 155.570 ;
        RECT 92.905 155.385 93.195 155.430 ;
        RECT 94.795 155.385 95.085 155.430 ;
        RECT 97.915 155.385 98.205 155.430 ;
        RECT 101.720 155.570 102.010 155.615 ;
        RECT 103.820 155.570 104.110 155.615 ;
        RECT 105.390 155.570 105.680 155.615 ;
        RECT 101.720 155.430 105.680 155.570 ;
        RECT 101.720 155.385 102.010 155.430 ;
        RECT 103.820 155.385 104.110 155.430 ;
        RECT 105.390 155.385 105.680 155.430 ;
        RECT 106.740 155.570 107.060 155.630 ;
        RECT 109.055 155.570 109.345 155.615 ;
        RECT 106.740 155.430 109.345 155.570 ;
        RECT 106.740 155.370 107.060 155.430 ;
        RECT 109.055 155.385 109.345 155.430 ;
        RECT 111.380 155.570 111.670 155.615 ;
        RECT 113.480 155.570 113.770 155.615 ;
        RECT 115.050 155.570 115.340 155.615 ;
        RECT 111.380 155.430 115.340 155.570 ;
        RECT 111.380 155.385 111.670 155.430 ;
        RECT 113.480 155.385 113.770 155.430 ;
        RECT 115.050 155.385 115.340 155.430 ;
        RECT 73.635 155.230 73.925 155.275 ;
        RECT 75.460 155.230 75.780 155.290 ;
        RECT 92.035 155.230 92.325 155.275 ;
        RECT 93.860 155.230 94.180 155.290 ;
        RECT 101.235 155.230 101.525 155.275 ;
        RECT 73.635 155.090 101.525 155.230 ;
        RECT 73.635 155.045 73.925 155.090 ;
        RECT 75.460 155.030 75.780 155.090 ;
        RECT 84.290 154.950 84.430 155.090 ;
        RECT 92.035 155.045 92.325 155.090 ;
        RECT 93.860 155.030 94.180 155.090 ;
        RECT 101.235 155.045 101.525 155.090 ;
        RECT 102.115 155.230 102.405 155.275 ;
        RECT 103.305 155.230 103.595 155.275 ;
        RECT 105.825 155.230 106.115 155.275 ;
        RECT 108.120 155.230 108.440 155.290 ;
        RECT 110.895 155.230 111.185 155.275 ;
        RECT 102.115 155.090 106.115 155.230 ;
        RECT 102.115 155.045 102.405 155.090 ;
        RECT 103.305 155.045 103.595 155.090 ;
        RECT 105.825 155.045 106.115 155.090 ;
        RECT 106.370 155.090 111.185 155.230 ;
        RECT 74.100 154.890 74.390 154.935 ;
        RECT 75.935 154.890 76.225 154.935 ;
        RECT 79.515 154.890 79.805 154.935 ;
        RECT 74.100 154.750 79.805 154.890 ;
        RECT 74.100 154.705 74.390 154.750 ;
        RECT 75.935 154.705 76.225 154.750 ;
        RECT 79.515 154.705 79.805 154.750 ;
        RECT 80.595 154.890 80.885 154.910 ;
        RECT 82.820 154.890 83.140 154.950 ;
        RECT 80.595 154.750 83.140 154.890 ;
        RECT 75.000 154.350 75.320 154.610 ;
        RECT 80.595 154.595 80.885 154.750 ;
        RECT 82.820 154.690 83.140 154.750 ;
        RECT 84.200 154.690 84.520 154.950 ;
        RECT 87.435 154.705 87.725 154.935 ;
        RECT 91.575 154.705 91.865 154.935 ;
        RECT 92.500 154.890 92.790 154.935 ;
        RECT 94.335 154.890 94.625 154.935 ;
        RECT 97.915 154.890 98.205 154.935 ;
        RECT 92.500 154.750 98.205 154.890 ;
        RECT 92.500 154.705 92.790 154.750 ;
        RECT 94.335 154.705 94.625 154.750 ;
        RECT 97.915 154.705 98.205 154.750 ;
        RECT 77.295 154.550 77.945 154.595 ;
        RECT 80.595 154.550 81.185 154.595 ;
        RECT 87.510 154.550 87.650 154.705 ;
        RECT 77.295 154.410 81.185 154.550 ;
        RECT 77.295 154.365 77.945 154.410 ;
        RECT 80.895 154.365 81.185 154.410 ;
        RECT 82.450 154.410 87.650 154.550 ;
        RECT 82.450 154.255 82.590 154.410 ;
        RECT 82.375 154.025 82.665 154.255 ;
        RECT 84.660 154.010 84.980 154.270 ;
        RECT 91.650 154.210 91.790 154.705 ;
        RECT 95.700 154.595 96.020 154.610 ;
        RECT 98.995 154.595 99.285 154.910 ;
        RECT 101.310 154.890 101.450 155.045 ;
        RECT 106.370 154.890 106.510 155.090 ;
        RECT 108.120 155.030 108.440 155.090 ;
        RECT 110.895 155.045 111.185 155.090 ;
        RECT 111.775 155.230 112.065 155.275 ;
        RECT 112.965 155.230 113.255 155.275 ;
        RECT 115.485 155.230 115.775 155.275 ;
        RECT 111.775 155.090 115.775 155.230 ;
        RECT 111.775 155.045 112.065 155.090 ;
        RECT 112.965 155.045 113.255 155.090 ;
        RECT 115.485 155.045 115.775 155.090 ;
        RECT 101.310 154.750 106.510 154.890 ;
        RECT 95.695 154.550 96.345 154.595 ;
        RECT 98.995 154.550 99.585 154.595 ;
        RECT 95.695 154.410 99.585 154.550 ;
        RECT 95.695 154.365 96.345 154.410 ;
        RECT 99.295 154.365 99.585 154.410 ;
        RECT 95.700 154.350 96.020 154.365 ;
        RECT 93.860 154.210 94.180 154.270 ;
        RECT 91.650 154.070 94.180 154.210 ;
        RECT 101.310 154.210 101.450 154.750 ;
        RECT 109.500 154.690 109.820 154.950 ;
        RECT 102.570 154.550 102.860 154.595 ;
        RECT 103.520 154.550 103.840 154.610 ;
        RECT 102.570 154.410 103.840 154.550 ;
        RECT 102.570 154.365 102.860 154.410 ;
        RECT 103.520 154.350 103.840 154.410 ;
        RECT 102.140 154.210 102.460 154.270 ;
        RECT 101.310 154.070 102.460 154.210 ;
        RECT 93.860 154.010 94.180 154.070 ;
        RECT 102.140 154.010 102.460 154.070 ;
        RECT 103.060 154.210 103.380 154.270 ;
        RECT 109.590 154.210 109.730 154.690 ;
        RECT 112.230 154.550 112.520 154.595 ;
        RECT 115.020 154.550 115.340 154.610 ;
        RECT 112.230 154.410 115.340 154.550 ;
        RECT 112.230 154.365 112.520 154.410 ;
        RECT 115.020 154.350 115.340 154.410 ;
        RECT 103.060 154.070 109.730 154.210 ;
        RECT 103.060 154.010 103.380 154.070 ;
        RECT 121.455 153.870 121.935 158.830 ;
        RECT 71.250 153.390 121.935 153.870 ;
        RECT 75.000 153.190 75.320 153.250 ;
        RECT 77.775 153.190 78.065 153.235 ;
        RECT 75.000 153.050 78.065 153.190 ;
        RECT 75.000 152.990 75.320 153.050 ;
        RECT 77.775 153.005 78.065 153.050 ;
        RECT 84.660 152.990 84.980 153.250 ;
        RECT 107.200 153.190 107.520 153.250 ;
        RECT 101.770 153.050 107.520 153.190 ;
        RECT 83.295 152.510 83.585 152.555 ;
        RECT 84.750 152.510 84.890 152.990 ;
        RECT 96.620 152.650 96.940 152.910 ;
        RECT 101.770 152.555 101.910 153.050 ;
        RECT 107.200 152.990 107.520 153.050 ;
        RECT 110.880 152.990 111.200 153.250 ;
        RECT 115.020 152.990 115.340 153.250 ;
        RECT 116.875 153.190 117.165 153.235 ;
        RECT 119.160 153.190 119.480 153.250 ;
        RECT 116.875 153.050 119.480 153.190 ;
        RECT 116.875 153.005 117.165 153.050 ;
        RECT 119.160 152.990 119.480 153.050 ;
        RECT 120.080 152.990 120.400 153.250 ;
        RECT 102.140 152.650 102.460 152.910 ;
        RECT 103.535 152.850 103.825 152.895 ;
        RECT 103.535 152.710 112.030 152.850 ;
        RECT 103.535 152.665 103.825 152.710 ;
        RECT 83.295 152.370 84.890 152.510 ;
        RECT 83.295 152.325 83.585 152.370 ;
        RECT 101.235 152.325 101.525 152.555 ;
        RECT 101.695 152.325 101.985 152.555 ;
        RECT 80.535 152.170 80.825 152.215 ;
        RECT 81.440 152.170 81.760 152.230 ;
        RECT 80.535 152.030 81.760 152.170 ;
        RECT 80.535 151.985 80.825 152.030 ;
        RECT 81.440 151.970 81.760 152.030 ;
        RECT 83.755 152.170 84.045 152.215 ;
        RECT 93.860 152.170 94.180 152.230 ;
        RECT 83.755 152.030 94.180 152.170 ;
        RECT 83.755 151.985 84.045 152.030 ;
        RECT 93.860 151.970 94.180 152.030 ;
        RECT 82.820 151.830 83.140 151.890 ;
        RECT 86.040 151.830 86.360 151.890 ;
        RECT 82.820 151.690 86.360 151.830 ;
        RECT 82.820 151.630 83.140 151.690 ;
        RECT 86.040 151.630 86.360 151.690 ;
        RECT 84.200 151.490 84.520 151.550 ;
        RECT 89.275 151.490 89.565 151.535 ;
        RECT 84.200 151.350 89.565 151.490 ;
        RECT 101.310 151.490 101.450 152.325 ;
        RECT 102.230 152.170 102.370 152.650 ;
        RECT 102.615 152.510 102.905 152.555 ;
        RECT 103.060 152.510 103.380 152.570 ;
        RECT 105.360 152.555 105.680 152.570 ;
        RECT 111.890 152.555 112.030 152.710 ;
        RECT 102.615 152.370 103.380 152.510 ;
        RECT 102.615 152.325 102.905 152.370 ;
        RECT 103.060 152.310 103.380 152.370 ;
        RECT 105.330 152.325 105.680 152.555 ;
        RECT 111.815 152.325 112.105 152.555 ;
        RECT 117.795 152.510 118.085 152.555 ;
        RECT 120.170 152.510 120.310 152.990 ;
        RECT 117.795 152.370 120.310 152.510 ;
        RECT 117.795 152.325 118.085 152.370 ;
        RECT 105.360 152.310 105.680 152.325 ;
        RECT 103.995 152.170 104.285 152.215 ;
        RECT 102.230 152.030 104.285 152.170 ;
        RECT 103.995 151.985 104.285 152.030 ;
        RECT 104.875 152.170 105.165 152.215 ;
        RECT 106.065 152.170 106.355 152.215 ;
        RECT 108.585 152.170 108.875 152.215 ;
        RECT 104.875 152.030 108.875 152.170 ;
        RECT 104.875 151.985 105.165 152.030 ;
        RECT 106.065 151.985 106.355 152.030 ;
        RECT 108.585 151.985 108.875 152.030 ;
        RECT 102.155 151.830 102.445 151.875 ;
        RECT 102.600 151.830 102.920 151.890 ;
        RECT 102.155 151.690 102.920 151.830 ;
        RECT 102.155 151.645 102.445 151.690 ;
        RECT 102.600 151.630 102.920 151.690 ;
        RECT 104.480 151.830 104.770 151.875 ;
        RECT 106.580 151.830 106.870 151.875 ;
        RECT 108.150 151.830 108.440 151.875 ;
        RECT 104.480 151.690 108.440 151.830 ;
        RECT 104.480 151.645 104.770 151.690 ;
        RECT 106.580 151.645 106.870 151.690 ;
        RECT 108.150 151.645 108.440 151.690 ;
        RECT 114.560 151.490 114.880 151.550 ;
        RECT 101.310 151.350 114.880 151.490 ;
        RECT 84.200 151.290 84.520 151.350 ;
        RECT 89.275 151.305 89.565 151.350 ;
        RECT 114.560 151.290 114.880 151.350 ;
        RECT 68.930 150.670 119.550 151.150 ;
        RECT 80.995 150.470 81.285 150.515 ;
        RECT 81.900 150.470 82.220 150.530 ;
        RECT 80.995 150.330 82.220 150.470 ;
        RECT 80.995 150.285 81.285 150.330 ;
        RECT 81.900 150.270 82.220 150.330 ;
        RECT 93.415 150.470 93.705 150.515 ;
        RECT 93.860 150.470 94.180 150.530 ;
        RECT 93.415 150.330 94.180 150.470 ;
        RECT 93.415 150.285 93.705 150.330 ;
        RECT 93.860 150.270 94.180 150.330 ;
        RECT 102.600 150.270 102.920 150.530 ;
        RECT 105.360 150.470 105.680 150.530 ;
        RECT 105.835 150.470 106.125 150.515 ;
        RECT 105.360 150.330 106.125 150.470 ;
        RECT 105.360 150.270 105.680 150.330 ;
        RECT 105.835 150.285 106.125 150.330 ;
        RECT 114.560 150.270 114.880 150.530 ;
        RECT 85.545 150.130 85.835 150.175 ;
        RECT 87.435 150.130 87.725 150.175 ;
        RECT 90.555 150.130 90.845 150.175 ;
        RECT 85.545 149.990 90.845 150.130 ;
        RECT 85.545 149.945 85.835 149.990 ;
        RECT 87.435 149.945 87.725 149.990 ;
        RECT 90.555 149.945 90.845 149.990 ;
        RECT 84.200 149.790 84.520 149.850 ;
        RECT 84.675 149.790 84.965 149.835 ;
        RECT 84.200 149.650 84.965 149.790 ;
        RECT 102.690 149.790 102.830 150.270 ;
        RECT 107.200 150.130 107.520 150.190 ;
        RECT 107.675 150.130 107.965 150.175 ;
        RECT 107.200 149.990 107.965 150.130 ;
        RECT 107.200 149.930 107.520 149.990 ;
        RECT 107.675 149.945 107.965 149.990 ;
        RECT 110.880 149.790 111.200 149.850 ;
        RECT 113.195 149.790 113.485 149.835 ;
        RECT 102.690 149.650 107.430 149.790 ;
        RECT 84.200 149.590 84.520 149.650 ;
        RECT 84.675 149.605 84.965 149.650 ;
        RECT 81.900 149.250 82.220 149.510 ;
        RECT 85.140 149.450 85.430 149.495 ;
        RECT 86.975 149.450 87.265 149.495 ;
        RECT 90.555 149.450 90.845 149.495 ;
        RECT 85.140 149.310 90.845 149.450 ;
        RECT 85.140 149.265 85.430 149.310 ;
        RECT 86.975 149.265 87.265 149.310 ;
        RECT 90.555 149.265 90.845 149.310 ;
        RECT 85.580 149.110 85.900 149.170 ;
        RECT 86.055 149.110 86.345 149.155 ;
        RECT 85.580 148.970 86.345 149.110 ;
        RECT 85.580 148.910 85.900 148.970 ;
        RECT 86.055 148.925 86.345 148.970 ;
        RECT 87.420 149.110 87.740 149.170 ;
        RECT 91.635 149.155 91.925 149.470 ;
        RECT 104.455 149.265 104.745 149.495 ;
        RECT 88.335 149.110 88.985 149.155 ;
        RECT 91.635 149.110 92.225 149.155 ;
        RECT 87.420 148.970 92.225 149.110 ;
        RECT 104.530 149.110 104.670 149.265 ;
        RECT 106.740 149.250 107.060 149.510 ;
        RECT 107.290 149.495 107.430 149.650 ;
        RECT 110.880 149.650 113.485 149.790 ;
        RECT 110.880 149.590 111.200 149.650 ;
        RECT 113.195 149.605 113.485 149.650 ;
        RECT 117.780 149.590 118.100 149.850 ;
        RECT 107.215 149.265 107.505 149.495 ;
        RECT 108.135 149.450 108.425 149.495 ;
        RECT 110.435 149.450 110.725 149.495 ;
        RECT 108.135 149.310 110.725 149.450 ;
        RECT 108.135 149.265 108.425 149.310 ;
        RECT 110.435 149.265 110.725 149.310 ;
        RECT 109.500 149.110 109.820 149.170 ;
        RECT 104.530 148.970 109.820 149.110 ;
        RECT 87.420 148.910 87.740 148.970 ;
        RECT 88.335 148.925 88.985 148.970 ;
        RECT 91.935 148.925 92.225 148.970 ;
        RECT 109.500 148.910 109.820 148.970 ;
        RECT 105.375 148.770 105.665 148.815 ;
        RECT 109.040 148.770 109.360 148.830 ;
        RECT 49.000 148.430 50.500 148.755 ;
        RECT 105.375 148.630 109.360 148.770 ;
        RECT 105.375 148.585 105.665 148.630 ;
        RECT 109.040 148.570 109.360 148.630 ;
        RECT 121.455 148.430 121.935 153.390 ;
        RECT 49.000 147.950 121.935 148.430 ;
        RECT 49.000 147.760 50.500 147.950 ;
        RECT 25.335 144.220 26.440 144.355 ;
        RECT 22.295 143.580 26.440 144.220 ;
        RECT 21.090 142.970 21.350 143.290 ;
        RECT 19.840 140.395 20.120 140.735 ;
        RECT 18.915 139.125 19.175 139.445 ;
        RECT 21.135 136.915 21.305 142.970 ;
        RECT 22.300 138.935 22.470 143.580 ;
        RECT 25.335 143.245 26.440 143.580 ;
        RECT 22.300 138.765 29.505 138.935 ;
        RECT 21.135 136.745 28.295 136.915 ;
        RECT 12.625 135.520 12.855 136.520 ;
        RECT 13.065 135.520 13.295 136.520 ;
        RECT 17.150 136.410 17.440 136.640 ;
        RECT 20.585 135.870 23.295 136.140 ;
        RECT 12.655 134.650 12.825 135.520 ;
        RECT 17.920 135.425 18.250 135.725 ;
        RECT 19.950 135.425 20.280 135.725 ;
        RECT 17.750 134.755 17.980 135.285 ;
        RECT 12.620 132.545 12.870 134.650 ;
        RECT 16.220 134.590 17.980 134.755 ;
        RECT 12.620 130.135 12.870 131.995 ;
        RECT 16.220 130.135 16.385 134.590 ;
        RECT 17.750 134.285 17.980 134.590 ;
        RECT 18.190 134.285 18.420 135.285 ;
        RECT 19.780 134.285 20.010 135.285 ;
        RECT 20.220 134.855 20.450 135.285 ;
        RECT 20.620 134.855 20.820 135.870 ;
        RECT 21.320 135.295 21.640 135.555 ;
        RECT 21.980 135.425 22.300 135.715 ;
        RECT 20.220 134.655 20.820 134.855 ;
        RECT 21.365 134.925 21.595 135.295 ;
        RECT 21.810 134.925 22.040 135.285 ;
        RECT 21.365 134.695 22.040 134.925 ;
        RECT 20.220 134.285 20.450 134.655 ;
        RECT 21.810 134.285 22.040 134.695 ;
        RECT 22.250 134.925 22.480 135.285 ;
        RECT 23.025 134.925 23.295 135.870 ;
        RECT 24.020 135.445 24.340 135.735 ;
        RECT 24.500 135.295 24.780 135.695 ;
        RECT 23.840 134.925 24.070 135.295 ;
        RECT 22.250 134.655 24.070 134.925 ;
        RECT 22.250 134.285 22.480 134.655 ;
        RECT 23.840 134.295 24.070 134.655 ;
        RECT 24.280 134.705 24.780 135.295 ;
        RECT 25.700 135.295 25.870 136.745 ;
        RECT 28.125 135.715 28.295 136.745 ;
        RECT 26.040 135.435 26.360 135.705 ;
        RECT 28.060 135.435 28.380 135.715 ;
        RECT 25.700 134.745 26.090 135.295 ;
        RECT 24.280 134.295 24.510 134.705 ;
        RECT 25.860 134.295 26.090 134.745 ;
        RECT 26.300 134.295 26.530 135.295 ;
        RECT 27.885 134.290 28.115 135.290 ;
        RECT 28.325 135.150 28.555 135.290 ;
        RECT 29.335 135.150 29.505 138.765 ;
        RECT 28.325 134.980 29.505 135.150 ;
        RECT 28.325 134.290 28.555 134.980 ;
        RECT 17.795 134.145 17.960 134.285 ;
        RECT 17.795 134.090 18.250 134.145 ;
        RECT 19.950 134.090 20.280 134.145 ;
        RECT 17.795 133.925 20.280 134.090 ;
        RECT 17.920 133.845 18.250 133.925 ;
        RECT 19.950 133.845 20.280 133.925 ;
        RECT 20.055 133.540 20.220 133.845 ;
        RECT 21.950 133.825 22.340 134.145 ;
        RECT 24.000 133.845 24.340 134.145 ;
        RECT 26.040 133.875 26.360 134.155 ;
        RECT 26.135 133.540 26.300 133.875 ;
        RECT 28.070 133.865 28.370 134.145 ;
        RECT 20.055 133.375 26.300 133.540 ;
        RECT 17.500 131.290 18.040 131.560 ;
        RECT 19.610 131.290 19.930 131.335 ;
        RECT 17.500 131.120 19.930 131.290 ;
        RECT 17.500 131.110 18.040 131.120 ;
        RECT 19.610 131.075 19.930 131.120 ;
        RECT 23.900 130.675 24.305 130.775 ;
        RECT 12.620 129.955 16.385 130.135 ;
        RECT 20.510 130.405 24.305 130.675 ;
        RECT 12.620 129.950 16.380 129.955 ;
        RECT 12.620 129.890 12.870 129.950 ;
        RECT 12.350 124.405 14.535 125.235 ;
        RECT 10.665 124.235 14.535 124.405 ;
        RECT 10.665 104.265 10.835 124.235 ;
        RECT 12.350 123.435 14.535 124.235 ;
        RECT 20.510 119.825 20.780 130.405 ;
        RECT 20.510 119.555 42.415 119.825 ;
        RECT 17.390 114.950 17.765 115.295 ;
        RECT 20.410 115.235 20.745 115.315 ;
        RECT 19.590 115.035 20.745 115.235 ;
        RECT 17.475 112.765 17.665 114.950 ;
        RECT 18.710 113.195 18.940 114.195 ;
        RECT 19.150 113.195 19.380 114.195 ;
        RECT 19.590 113.195 19.820 115.035 ;
        RECT 20.410 114.970 20.745 115.035 ;
        RECT 20.220 113.195 20.450 114.195 ;
        RECT 20.660 113.195 20.890 114.195 ;
        RECT 21.100 113.490 21.330 114.195 ;
        RECT 21.100 113.320 22.250 113.490 ;
        RECT 21.100 113.195 21.330 113.320 ;
        RECT 18.740 112.765 18.910 113.195 ;
        RECT 17.475 112.600 18.920 112.765 ;
        RECT 14.230 108.720 15.745 109.985 ;
        RECT 10.665 104.095 17.160 104.265 ;
        RECT 16.990 98.670 17.160 104.095 ;
        RECT 18.740 101.475 18.910 112.600 ;
        RECT 19.620 109.955 19.790 113.195 ;
        RECT 20.250 112.520 20.420 113.195 ;
        RECT 20.880 112.520 21.110 112.580 ;
        RECT 20.250 112.350 21.110 112.520 ;
        RECT 20.250 112.165 20.420 112.350 ;
        RECT 20.880 112.290 21.110 112.350 ;
        RECT 20.205 111.845 20.465 112.165 ;
        RECT 19.380 109.535 19.830 109.955 ;
        RECT 19.620 102.765 19.790 109.535 ;
        RECT 22.080 106.250 22.250 113.320 ;
        RECT 25.115 106.250 26.220 106.385 ;
        RECT 22.075 105.610 26.220 106.250 ;
        RECT 20.870 105.000 21.130 105.320 ;
        RECT 19.620 102.425 19.900 102.765 ;
        RECT 18.695 101.155 18.955 101.475 ;
        RECT 20.915 98.945 21.085 105.000 ;
        RECT 22.080 100.965 22.250 105.610 ;
        RECT 25.115 105.275 26.220 105.610 ;
        RECT 22.080 100.795 29.285 100.965 ;
        RECT 20.915 98.775 28.075 98.945 ;
        RECT 12.405 97.550 12.635 98.550 ;
        RECT 12.845 97.550 13.075 98.550 ;
        RECT 16.930 98.440 17.220 98.670 ;
        RECT 20.365 97.900 23.075 98.170 ;
        RECT 12.435 96.680 12.605 97.550 ;
        RECT 17.700 97.455 18.030 97.755 ;
        RECT 19.730 97.455 20.060 97.755 ;
        RECT 17.530 96.785 17.760 97.315 ;
        RECT 12.400 94.575 12.650 96.680 ;
        RECT 16.000 96.620 17.760 96.785 ;
        RECT 12.400 92.165 12.650 94.025 ;
        RECT 16.000 92.165 16.165 96.620 ;
        RECT 17.530 96.315 17.760 96.620 ;
        RECT 17.970 96.315 18.200 97.315 ;
        RECT 19.560 96.315 19.790 97.315 ;
        RECT 20.000 96.885 20.230 97.315 ;
        RECT 20.400 96.885 20.600 97.900 ;
        RECT 21.100 97.325 21.420 97.585 ;
        RECT 21.760 97.455 22.080 97.745 ;
        RECT 20.000 96.685 20.600 96.885 ;
        RECT 21.145 96.955 21.375 97.325 ;
        RECT 21.590 96.955 21.820 97.315 ;
        RECT 21.145 96.725 21.820 96.955 ;
        RECT 20.000 96.315 20.230 96.685 ;
        RECT 21.590 96.315 21.820 96.725 ;
        RECT 22.030 96.955 22.260 97.315 ;
        RECT 22.805 96.955 23.075 97.900 ;
        RECT 23.800 97.475 24.120 97.765 ;
        RECT 24.280 97.325 24.560 97.725 ;
        RECT 23.620 96.955 23.850 97.325 ;
        RECT 22.030 96.685 23.850 96.955 ;
        RECT 22.030 96.315 22.260 96.685 ;
        RECT 23.620 96.325 23.850 96.685 ;
        RECT 24.060 96.735 24.560 97.325 ;
        RECT 25.480 97.325 25.650 98.775 ;
        RECT 27.905 97.745 28.075 98.775 ;
        RECT 25.820 97.465 26.140 97.735 ;
        RECT 27.840 97.465 28.160 97.745 ;
        RECT 25.480 96.775 25.870 97.325 ;
        RECT 24.060 96.325 24.290 96.735 ;
        RECT 25.640 96.325 25.870 96.775 ;
        RECT 26.080 96.325 26.310 97.325 ;
        RECT 27.665 96.320 27.895 97.320 ;
        RECT 28.105 97.180 28.335 97.320 ;
        RECT 29.115 97.180 29.285 100.795 ;
        RECT 28.105 97.010 29.285 97.180 ;
        RECT 28.105 96.320 28.335 97.010 ;
        RECT 17.575 96.175 17.740 96.315 ;
        RECT 17.575 96.120 18.030 96.175 ;
        RECT 19.730 96.120 20.060 96.175 ;
        RECT 17.575 95.955 20.060 96.120 ;
        RECT 17.700 95.875 18.030 95.955 ;
        RECT 19.730 95.875 20.060 95.955 ;
        RECT 19.835 95.570 20.000 95.875 ;
        RECT 21.730 95.855 22.120 96.175 ;
        RECT 23.780 95.875 24.120 96.175 ;
        RECT 25.820 95.905 26.140 96.185 ;
        RECT 25.915 95.570 26.080 95.905 ;
        RECT 27.850 95.895 28.150 96.175 ;
        RECT 19.835 95.405 26.080 95.570 ;
        RECT 17.400 93.320 17.570 93.555 ;
        RECT 19.390 93.320 19.710 93.365 ;
        RECT 17.400 93.150 19.710 93.320 ;
        RECT 17.400 93.145 17.570 93.150 ;
        RECT 19.390 93.105 19.710 93.150 ;
        RECT 23.680 92.705 24.085 92.805 ;
        RECT 12.400 91.985 16.165 92.165 ;
        RECT 20.290 92.435 24.085 92.705 ;
        RECT 12.400 91.980 16.160 91.985 ;
        RECT 12.400 91.920 12.650 91.980 ;
        RECT 1.000 83.125 2.500 83.410 ;
        RECT 20.290 83.125 20.560 92.435 ;
        RECT 42.145 83.125 42.415 119.555 ;
        RECT 49.000 89.180 50.500 89.630 ;
        RECT 49.000 88.700 152.240 89.180 ;
        RECT 49.000 88.690 89.620 88.700 ;
        RECT 49.000 88.350 50.500 88.690 ;
        RECT 88.980 83.740 89.460 88.690 ;
        RECT 103.550 88.500 103.870 88.560 ;
        RECT 104.945 88.500 105.235 88.545 ;
        RECT 103.550 88.360 105.235 88.500 ;
        RECT 103.550 88.300 103.870 88.360 ;
        RECT 104.945 88.315 105.235 88.360 ;
        RECT 139.430 88.500 139.750 88.560 ;
        RECT 140.825 88.500 141.115 88.545 ;
        RECT 139.430 88.360 141.115 88.500 ;
        RECT 139.430 88.300 139.750 88.360 ;
        RECT 140.825 88.315 141.115 88.360 ;
        RECT 150.025 88.160 150.315 88.205 ;
        RECT 151.850 88.160 152.170 88.220 ;
        RECT 150.025 88.020 152.170 88.160 ;
        RECT 150.025 87.975 150.315 88.020 ;
        RECT 151.850 87.960 152.170 88.020 ;
        RECT 106.310 87.620 106.630 87.880 ;
        RECT 140.350 87.620 140.670 87.880 ;
        RECT 145.870 87.140 146.190 87.200 ;
        RECT 149.105 87.140 149.395 87.185 ;
        RECT 145.870 87.000 149.395 87.140 ;
        RECT 145.870 86.940 146.190 87.000 ;
        RECT 149.105 86.955 149.395 87.000 ;
        RECT 91.060 85.980 153.380 86.460 ;
        RECT 137.555 85.440 137.845 85.485 ;
        RECT 139.445 85.440 139.735 85.485 ;
        RECT 142.565 85.440 142.855 85.485 ;
        RECT 137.555 85.300 142.855 85.440 ;
        RECT 137.555 85.255 137.845 85.300 ;
        RECT 139.445 85.255 139.735 85.300 ;
        RECT 142.565 85.255 142.855 85.300 ;
        RECT 118.270 85.100 118.590 85.160 ;
        RECT 125.630 85.100 125.950 85.160 ;
        RECT 136.685 85.100 136.975 85.145 ;
        RECT 118.270 84.960 120.110 85.100 ;
        RECT 118.270 84.900 118.590 84.960 ;
        RECT 119.970 84.420 120.110 84.960 ;
        RECT 125.630 84.960 136.975 85.100 ;
        RECT 125.630 84.900 125.950 84.960 ;
        RECT 136.685 84.915 136.975 84.960 ;
        RECT 121.950 84.560 122.270 84.820 ;
        RECT 122.410 84.760 122.730 84.820 ;
        RECT 122.885 84.760 123.175 84.805 ;
        RECT 122.410 84.620 123.175 84.760 ;
        RECT 122.410 84.560 122.730 84.620 ;
        RECT 122.885 84.575 123.175 84.620 ;
        RECT 126.090 84.560 126.410 84.820 ;
        RECT 130.245 84.575 130.535 84.805 ;
        RECT 131.165 84.575 131.455 84.805 ;
        RECT 132.085 84.760 132.375 84.805 ;
        RECT 133.925 84.760 134.215 84.805 ;
        RECT 132.085 84.620 134.215 84.760 ;
        RECT 132.085 84.575 132.375 84.620 ;
        RECT 133.925 84.575 134.215 84.620 ;
        RECT 137.150 84.760 137.440 84.805 ;
        RECT 138.985 84.760 139.275 84.805 ;
        RECT 142.565 84.760 142.855 84.805 ;
        RECT 137.150 84.620 142.855 84.760 ;
        RECT 137.150 84.575 137.440 84.620 ;
        RECT 138.985 84.575 139.275 84.620 ;
        RECT 142.565 84.575 142.855 84.620 ;
        RECT 143.570 84.780 143.890 84.820 ;
        RECT 130.320 84.420 130.460 84.575 ;
        RECT 119.970 84.280 130.460 84.420 ;
        RECT 122.870 83.880 123.190 84.140 ;
        RECT 124.710 84.080 125.030 84.140 ;
        RECT 125.185 84.080 125.475 84.125 ;
        RECT 124.710 83.940 125.475 84.080 ;
        RECT 124.710 83.880 125.030 83.940 ;
        RECT 125.185 83.895 125.475 83.940 ;
        RECT 127.470 84.080 127.790 84.140 ;
        RECT 131.240 84.080 131.380 84.575 ;
        RECT 143.570 84.560 143.935 84.780 ;
        RECT 143.645 84.465 143.935 84.560 ;
        RECT 138.065 84.235 138.355 84.465 ;
        RECT 140.345 84.420 140.995 84.465 ;
        RECT 143.645 84.420 144.235 84.465 ;
        RECT 140.345 84.280 144.235 84.420 ;
        RECT 140.345 84.235 140.995 84.280 ;
        RECT 143.945 84.235 144.235 84.280 ;
        RECT 127.470 83.940 131.380 84.080 ;
        RECT 134.845 84.080 135.135 84.125 ;
        RECT 138.140 84.080 138.280 84.235 ;
        RECT 134.845 83.940 138.280 84.080 ;
        RECT 127.470 83.880 127.790 83.940 ;
        RECT 134.845 83.895 135.135 83.940 ;
        RECT 145.410 83.880 145.730 84.140 ;
        RECT 88.980 83.260 152.240 83.740 ;
        RECT 1.000 82.855 42.445 83.125 ;
        RECT 1.000 82.850 20.495 82.855 ;
        RECT 1.000 82.525 2.500 82.850 ;
        RECT 88.980 78.300 89.460 83.260 ;
        RECT 122.410 83.060 122.730 83.120 ;
        RECT 122.410 82.920 131.840 83.060 ;
        RECT 122.410 82.860 122.730 82.920 ;
        RECT 118.205 82.720 118.495 82.765 ;
        RECT 118.730 82.720 119.050 82.780 ;
        RECT 118.205 82.580 119.050 82.720 ;
        RECT 118.205 82.535 118.495 82.580 ;
        RECT 118.730 82.520 119.050 82.580 ;
        RECT 119.205 82.535 119.495 82.765 ;
        RECT 120.585 82.720 120.875 82.765 ;
        RECT 121.950 82.720 122.270 82.780 ;
        RECT 120.585 82.580 122.270 82.720 ;
        RECT 120.585 82.535 120.875 82.580 ;
        RECT 113.685 82.195 113.975 82.425 ;
        RECT 115.985 82.380 116.275 82.425 ;
        RECT 115.985 82.240 117.580 82.380 ;
        RECT 115.985 82.195 116.275 82.240 ;
        RECT 113.210 82.040 113.530 82.100 ;
        RECT 113.760 82.040 113.900 82.195 ;
        RECT 113.210 81.900 113.900 82.040 ;
        RECT 114.145 82.040 114.435 82.085 ;
        RECT 115.050 82.040 115.370 82.100 ;
        RECT 114.145 81.900 115.370 82.040 ;
        RECT 113.210 81.840 113.530 81.900 ;
        RECT 114.145 81.855 114.435 81.900 ;
        RECT 115.050 81.840 115.370 81.900 ;
        RECT 117.440 81.745 117.580 82.240 ;
        RECT 118.270 82.040 118.590 82.100 ;
        RECT 119.280 82.040 119.420 82.535 ;
        RECT 121.950 82.520 122.270 82.580 ;
        RECT 121.505 82.380 121.795 82.425 ;
        RECT 122.500 82.380 122.640 82.860 ;
        RECT 125.630 82.720 125.950 82.780 ;
        RECT 122.960 82.580 125.950 82.720 ;
        RECT 122.960 82.425 123.100 82.580 ;
        RECT 125.630 82.520 125.950 82.580 ;
        RECT 126.545 82.720 127.195 82.765 ;
        RECT 127.930 82.720 128.250 82.780 ;
        RECT 130.145 82.720 130.435 82.765 ;
        RECT 126.545 82.580 130.435 82.720 ;
        RECT 126.545 82.535 127.195 82.580 ;
        RECT 127.930 82.520 128.250 82.580 ;
        RECT 129.845 82.535 130.435 82.580 ;
        RECT 121.505 82.240 122.640 82.380 ;
        RECT 121.505 82.195 121.795 82.240 ;
        RECT 122.885 82.195 123.175 82.425 ;
        RECT 123.350 82.380 123.640 82.425 ;
        RECT 125.185 82.380 125.475 82.425 ;
        RECT 128.765 82.380 129.055 82.425 ;
        RECT 123.350 82.240 129.055 82.380 ;
        RECT 123.350 82.195 123.640 82.240 ;
        RECT 125.185 82.195 125.475 82.240 ;
        RECT 128.765 82.195 129.055 82.240 ;
        RECT 129.845 82.220 130.135 82.535 ;
        RECT 118.270 81.900 119.420 82.040 ;
        RECT 124.265 82.040 124.555 82.085 ;
        RECT 124.710 82.040 125.030 82.100 ;
        RECT 131.700 82.085 131.840 82.920 ;
        RECT 143.570 82.860 143.890 83.120 ;
        RECT 139.060 82.580 146.100 82.720 ;
        RECT 133.910 82.380 134.230 82.440 ;
        RECT 139.060 82.425 139.200 82.580 ;
        RECT 145.960 82.440 146.100 82.580 ;
        RECT 134.385 82.380 134.675 82.425 ;
        RECT 133.910 82.240 134.675 82.380 ;
        RECT 133.910 82.180 134.230 82.240 ;
        RECT 134.385 82.195 134.675 82.240 ;
        RECT 138.985 82.195 139.275 82.425 ;
        RECT 142.650 82.380 142.970 82.440 ;
        RECT 144.045 82.380 144.335 82.425 ;
        RECT 142.650 82.240 144.335 82.380 ;
        RECT 142.650 82.180 142.970 82.240 ;
        RECT 144.045 82.195 144.335 82.240 ;
        RECT 145.870 82.180 146.190 82.440 ;
        RECT 124.265 81.900 125.030 82.040 ;
        RECT 118.270 81.840 118.590 81.900 ;
        RECT 124.265 81.855 124.555 81.900 ;
        RECT 124.710 81.840 125.030 81.900 ;
        RECT 131.625 82.040 131.915 82.085 ;
        RECT 133.005 82.040 133.295 82.085 ;
        RECT 136.210 82.040 136.530 82.100 ;
        RECT 131.625 81.900 136.530 82.040 ;
        RECT 131.625 81.855 131.915 81.900 ;
        RECT 133.005 81.855 133.295 81.900 ;
        RECT 136.210 81.840 136.530 81.900 ;
        RECT 117.365 81.515 117.655 81.745 ;
        RECT 123.755 81.700 124.045 81.745 ;
        RECT 125.645 81.700 125.935 81.745 ;
        RECT 128.765 81.700 129.055 81.745 ;
        RECT 123.755 81.560 129.055 81.700 ;
        RECT 123.755 81.515 124.045 81.560 ;
        RECT 125.645 81.515 125.935 81.560 ;
        RECT 128.765 81.515 129.055 81.560 ;
        RECT 133.465 81.700 133.755 81.745 ;
        RECT 134.830 81.700 135.150 81.760 ;
        RECT 138.525 81.700 138.815 81.745 ;
        RECT 133.465 81.560 138.815 81.700 ;
        RECT 133.465 81.515 133.755 81.560 ;
        RECT 134.830 81.500 135.150 81.560 ;
        RECT 138.525 81.515 138.815 81.560 ;
        RECT 115.065 81.360 115.355 81.405 ;
        RECT 115.510 81.360 115.830 81.420 ;
        RECT 115.065 81.220 115.830 81.360 ;
        RECT 115.065 81.175 115.355 81.220 ;
        RECT 115.510 81.160 115.830 81.220 ;
        RECT 118.285 81.360 118.575 81.405 ;
        RECT 121.490 81.360 121.810 81.420 ;
        RECT 118.285 81.220 121.810 81.360 ;
        RECT 118.285 81.175 118.575 81.220 ;
        RECT 121.490 81.160 121.810 81.220 ;
        RECT 122.410 81.160 122.730 81.420 ;
        RECT 135.305 81.360 135.595 81.405 ;
        RECT 137.130 81.360 137.450 81.420 ;
        RECT 135.305 81.220 137.450 81.360 ;
        RECT 135.305 81.175 135.595 81.220 ;
        RECT 137.130 81.160 137.450 81.220 ;
        RECT 152.900 81.020 153.380 85.980 ;
        RECT 91.060 80.540 153.380 81.020 ;
        RECT 122.425 80.340 122.715 80.385 ;
        RECT 122.870 80.340 123.190 80.400 ;
        RECT 127.930 80.340 128.250 80.400 ;
        RECT 128.405 80.340 128.695 80.385 ;
        RECT 122.425 80.200 126.320 80.340 ;
        RECT 122.425 80.155 122.715 80.200 ;
        RECT 122.870 80.140 123.190 80.200 ;
        RECT 111.795 80.000 112.085 80.045 ;
        RECT 113.685 80.000 113.975 80.045 ;
        RECT 116.805 80.000 117.095 80.045 ;
        RECT 111.795 79.860 117.095 80.000 ;
        RECT 111.795 79.815 112.085 79.860 ;
        RECT 113.685 79.815 113.975 79.860 ;
        RECT 116.805 79.815 117.095 79.860 ;
        RECT 117.900 79.860 123.100 80.000 ;
        RECT 110.910 79.660 111.230 79.720 ;
        RECT 117.900 79.660 118.040 79.860 ;
        RECT 110.910 79.520 118.040 79.660 ;
        RECT 110.910 79.460 111.230 79.520 ;
        RECT 118.270 79.460 118.590 79.720 ;
        RECT 111.390 79.320 111.680 79.365 ;
        RECT 113.225 79.320 113.515 79.365 ;
        RECT 116.805 79.320 117.095 79.365 ;
        RECT 111.390 79.180 117.095 79.320 ;
        RECT 111.390 79.135 111.680 79.180 ;
        RECT 113.225 79.135 113.515 79.180 ;
        RECT 116.805 79.135 117.095 79.180 ;
        RECT 115.050 79.025 115.370 79.040 ;
        RECT 112.305 78.795 112.595 79.025 ;
        RECT 114.585 78.980 115.370 79.025 ;
        RECT 117.885 79.025 118.175 79.340 ;
        RECT 118.360 79.320 118.500 79.460 ;
        RECT 119.190 79.320 119.510 79.380 ;
        RECT 122.960 79.320 123.100 79.860 ;
        RECT 123.345 79.815 123.635 80.045 ;
        RECT 123.420 79.660 123.560 79.815 ;
        RECT 126.180 79.705 126.320 80.200 ;
        RECT 127.930 80.200 128.695 80.340 ;
        RECT 127.930 80.140 128.250 80.200 ;
        RECT 128.405 80.155 128.695 80.200 ;
        RECT 133.910 80.140 134.230 80.400 ;
        RECT 137.590 80.340 137.910 80.400 ;
        RECT 134.460 80.200 137.910 80.340 ;
        RECT 127.470 79.800 127.790 80.060 ;
        RECT 134.460 80.045 134.600 80.200 ;
        RECT 137.590 80.140 137.910 80.200 ;
        RECT 144.965 80.340 145.255 80.385 ;
        RECT 145.410 80.340 145.730 80.400 ;
        RECT 144.965 80.200 145.730 80.340 ;
        RECT 144.965 80.155 145.255 80.200 ;
        RECT 134.385 79.815 134.675 80.045 ;
        RECT 145.040 80.000 145.180 80.155 ;
        RECT 145.410 80.140 145.730 80.200 ;
        RECT 134.920 79.860 145.180 80.000 ;
        RECT 123.420 79.520 124.940 79.660 ;
        RECT 124.250 79.320 124.570 79.380 ;
        RECT 118.360 79.180 121.720 79.320 ;
        RECT 122.960 79.180 124.570 79.320 ;
        RECT 119.190 79.120 119.510 79.180 ;
        RECT 121.580 79.025 121.720 79.180 ;
        RECT 124.250 79.120 124.570 79.180 ;
        RECT 122.410 79.025 122.730 79.040 ;
        RECT 117.885 78.980 118.475 79.025 ;
        RECT 114.585 78.840 118.475 78.980 ;
        RECT 114.585 78.795 115.370 78.840 ;
        RECT 118.185 78.795 118.475 78.840 ;
        RECT 121.505 78.795 121.795 79.025 ;
        RECT 122.410 78.795 122.795 79.025 ;
        RECT 124.800 78.980 124.940 79.520 ;
        RECT 126.105 79.475 126.395 79.705 ;
        RECT 134.920 79.660 135.060 79.860 ;
        RECT 127.560 79.520 135.060 79.660 ;
        RECT 125.645 79.320 125.935 79.365 ;
        RECT 127.560 79.320 127.700 79.520 ;
        RECT 125.645 79.180 127.700 79.320 ;
        RECT 125.645 79.135 125.935 79.180 ;
        RECT 127.945 79.135 128.235 79.365 ;
        RECT 126.090 78.980 126.410 79.040 ;
        RECT 124.800 78.840 126.410 78.980 ;
        RECT 112.380 78.640 112.520 78.795 ;
        RECT 115.050 78.780 115.370 78.795 ;
        RECT 122.410 78.780 122.730 78.795 ;
        RECT 126.090 78.780 126.410 78.840 ;
        RECT 127.470 78.980 127.790 79.040 ;
        RECT 128.020 78.980 128.160 79.135 ;
        RECT 131.150 79.120 131.470 79.380 ;
        RECT 133.005 79.135 133.295 79.365 ;
        RECT 134.830 79.320 135.150 79.380 ;
        RECT 136.210 79.365 136.530 79.380 ;
        RECT 137.195 79.370 137.485 79.415 ;
        RECT 137.680 79.370 137.820 79.860 ;
        RECT 135.305 79.320 135.595 79.365 ;
        RECT 134.830 79.180 135.595 79.320 ;
        RECT 127.470 78.840 128.160 78.980 ;
        RECT 130.690 78.980 131.010 79.040 ;
        RECT 132.085 78.980 132.375 79.025 ;
        RECT 130.690 78.840 132.375 78.980 ;
        RECT 127.470 78.780 127.790 78.840 ;
        RECT 130.690 78.780 131.010 78.840 ;
        RECT 132.085 78.795 132.375 78.840 ;
        RECT 132.545 78.795 132.835 79.025 ;
        RECT 133.080 78.980 133.220 79.135 ;
        RECT 134.830 79.120 135.150 79.180 ;
        RECT 135.305 79.135 135.595 79.180 ;
        RECT 136.130 79.135 136.530 79.365 ;
        RECT 136.685 79.135 136.975 79.365 ;
        RECT 137.195 79.230 137.820 79.370 ;
        RECT 145.425 79.320 145.715 79.365 ;
        RECT 145.870 79.320 146.190 79.380 ;
        RECT 137.195 79.185 137.485 79.230 ;
        RECT 145.425 79.180 146.190 79.320 ;
        RECT 145.425 79.135 145.715 79.180 ;
        RECT 136.210 79.120 136.530 79.135 ;
        RECT 133.080 78.840 135.520 78.980 ;
        RECT 115.510 78.640 115.830 78.700 ;
        RECT 112.380 78.500 115.830 78.640 ;
        RECT 115.510 78.440 115.830 78.500 ;
        RECT 119.665 78.640 119.955 78.685 ;
        RECT 121.030 78.640 121.350 78.700 ;
        RECT 132.620 78.640 132.760 78.795 ;
        RECT 135.380 78.700 135.520 78.840 ;
        RECT 133.680 78.640 134.000 78.700 ;
        RECT 119.665 78.500 134.000 78.640 ;
        RECT 119.665 78.455 119.955 78.500 ;
        RECT 121.030 78.440 121.350 78.500 ;
        RECT 133.680 78.440 134.000 78.500 ;
        RECT 135.290 78.440 135.610 78.700 ;
        RECT 136.760 78.640 136.900 79.135 ;
        RECT 145.870 79.120 146.190 79.180 ;
        RECT 137.130 78.640 137.450 78.700 ;
        RECT 136.760 78.500 137.450 78.640 ;
        RECT 137.130 78.440 137.450 78.500 ;
        RECT 143.110 78.440 143.430 78.700 ;
        RECT 88.980 77.820 152.240 78.300 ;
        RECT 7.390 72.950 8.255 73.120 ;
        RECT 7.390 72.780 35.720 72.950 ;
        RECT 7.390 72.580 8.255 72.780 ;
        RECT 23.400 71.850 23.830 72.300 ;
        RECT 32.795 71.800 33.470 72.475 ;
        RECT 21.860 69.350 22.090 70.350 ;
        RECT 22.300 69.350 22.530 70.350 ;
        RECT 24.280 69.630 24.510 70.630 ;
        RECT 24.720 69.630 24.950 70.630 ;
        RECT 25.160 69.630 25.390 70.630 ;
        RECT 7.400 68.840 8.250 69.155 ;
        RECT 26.150 68.940 26.380 69.940 ;
        RECT 26.590 68.940 26.820 69.940 ;
        RECT 27.400 69.580 28.085 70.140 ;
        RECT 29.610 69.630 29.840 70.630 ;
        RECT 30.050 69.630 30.280 70.630 ;
        RECT 30.490 69.630 30.720 70.630 ;
        RECT 34.260 70.370 34.630 70.450 ;
        RECT 31.165 70.225 34.630 70.370 ;
        RECT 31.165 69.495 31.310 70.225 ;
        RECT 34.260 70.140 34.630 70.225 ;
        RECT 31.035 69.155 31.405 69.495 ;
        RECT 31.720 68.940 31.950 69.940 ;
        RECT 32.160 68.940 32.390 69.940 ;
        RECT 32.770 68.940 33.000 69.940 ;
        RECT 33.210 68.940 33.440 69.940 ;
        RECT 7.400 68.595 20.380 68.840 ;
        RECT 7.400 68.395 8.250 68.595 ;
        RECT 20.135 67.310 20.380 68.595 ;
        RECT 21.860 67.680 22.090 68.680 ;
        RECT 22.300 67.680 22.530 68.680 ;
        RECT 24.280 67.680 24.510 68.680 ;
        RECT 24.720 67.680 24.950 68.680 ;
        RECT 25.160 67.680 25.390 68.680 ;
        RECT 19.990 66.940 20.500 67.310 ;
        RECT 26.150 67.270 26.380 68.270 ;
        RECT 26.590 67.270 26.820 68.270 ;
        RECT 27.310 67.270 27.900 67.900 ;
        RECT 29.610 67.680 29.840 68.680 ;
        RECT 30.050 67.680 30.280 68.680 ;
        RECT 30.490 67.680 30.720 68.680 ;
        RECT 31.720 67.270 31.950 68.270 ;
        RECT 32.160 67.270 32.390 68.270 ;
        RECT 32.770 67.270 33.000 68.270 ;
        RECT 33.210 67.270 33.440 68.270 ;
        RECT 31.665 66.885 32.005 66.935 ;
        RECT 33.840 66.905 34.250 66.985 ;
        RECT 35.550 66.905 35.720 72.780 ;
        RECT 33.840 66.885 35.720 66.905 ;
        RECT 31.665 66.735 35.720 66.885 ;
        RECT 88.980 72.860 89.460 77.820 ;
        RECT 118.820 77.480 120.340 77.620 ;
        RECT 118.820 77.325 118.960 77.480 ;
        RECT 118.745 77.095 119.035 77.325 ;
        RECT 119.745 77.280 120.035 77.325 ;
        RECT 119.280 77.140 120.035 77.280 ;
        RECT 109.545 76.940 109.835 76.985 ;
        RECT 115.050 76.940 115.370 77.000 ;
        RECT 109.545 76.800 115.370 76.940 ;
        RECT 109.545 76.755 109.835 76.800 ;
        RECT 115.050 76.740 115.370 76.800 ;
        RECT 118.270 76.940 118.590 77.000 ;
        RECT 119.280 76.940 119.420 77.140 ;
        RECT 119.745 77.095 120.035 77.140 ;
        RECT 118.270 76.800 119.420 76.940 ;
        RECT 120.200 76.940 120.340 77.480 ;
        RECT 120.585 77.435 120.875 77.665 ;
        RECT 120.660 77.280 120.800 77.435 ;
        RECT 121.490 77.420 121.810 77.680 ;
        RECT 121.950 77.420 122.270 77.680 ;
        RECT 132.990 77.420 133.310 77.680 ;
        RECT 135.750 77.620 136.070 77.680 ;
        RECT 134.920 77.480 136.070 77.620 ;
        RECT 122.040 77.280 122.180 77.420 ;
        RECT 120.660 77.140 122.180 77.280 ;
        RECT 121.030 76.940 121.350 77.000 ;
        RECT 122.040 76.985 122.180 77.140 ;
        RECT 133.080 76.985 133.220 77.420 ;
        RECT 134.385 77.280 134.675 77.325 ;
        RECT 134.920 77.280 135.060 77.480 ;
        RECT 135.750 77.420 136.070 77.480 ;
        RECT 136.670 77.620 136.990 77.680 ;
        RECT 136.670 77.480 141.040 77.620 ;
        RECT 136.670 77.420 136.990 77.480 ;
        RECT 134.385 77.140 135.060 77.280 ;
        RECT 137.220 77.140 140.580 77.280 ;
        RECT 134.385 77.095 134.675 77.140 ;
        RECT 120.200 76.800 121.350 76.940 ;
        RECT 118.270 76.740 118.590 76.800 ;
        RECT 121.030 76.740 121.350 76.800 ;
        RECT 121.965 76.755 122.255 76.985 ;
        RECT 132.545 76.755 132.835 76.985 ;
        RECT 133.005 76.755 133.295 76.985 ;
        RECT 113.210 76.600 113.530 76.660 ;
        RECT 127.470 76.600 127.790 76.660 ;
        RECT 113.210 76.460 127.790 76.600 ;
        RECT 113.210 76.400 113.530 76.460 ;
        RECT 127.470 76.400 127.790 76.460 ;
        RECT 131.150 76.400 131.470 76.660 ;
        RECT 132.620 76.600 132.760 76.755 ;
        RECT 133.450 76.740 133.770 77.000 ;
        RECT 135.290 76.940 135.610 77.000 ;
        RECT 135.765 76.940 136.055 76.985 ;
        RECT 135.290 76.800 136.055 76.940 ;
        RECT 135.290 76.740 135.610 76.800 ;
        RECT 135.765 76.755 136.055 76.800 ;
        RECT 136.210 76.940 136.530 77.000 ;
        RECT 137.220 76.940 137.360 77.140 ;
        RECT 140.440 77.000 140.580 77.140 ;
        RECT 136.210 76.800 137.360 76.940 ;
        RECT 135.840 76.600 135.980 76.755 ;
        RECT 136.210 76.740 136.530 76.800 ;
        RECT 137.590 76.740 137.910 77.000 ;
        RECT 140.350 76.740 140.670 77.000 ;
        RECT 140.900 76.985 141.040 77.480 ;
        RECT 145.410 77.420 145.730 77.680 ;
        RECT 140.825 76.940 141.115 76.985 ;
        RECT 144.045 76.940 144.335 76.985 ;
        RECT 140.825 76.800 144.335 76.940 ;
        RECT 145.500 76.940 145.640 77.420 ;
        RECT 146.345 76.940 146.635 76.985 ;
        RECT 145.500 76.800 146.635 76.940 ;
        RECT 140.825 76.755 141.115 76.800 ;
        RECT 144.045 76.755 144.335 76.800 ;
        RECT 146.345 76.755 146.635 76.800 ;
        RECT 142.205 76.600 142.495 76.645 ;
        RECT 143.110 76.600 143.430 76.660 ;
        RECT 132.620 76.460 133.220 76.600 ;
        RECT 131.240 76.260 131.380 76.400 ;
        RECT 133.080 76.260 133.220 76.460 ;
        RECT 135.840 76.460 141.500 76.600 ;
        RECT 135.840 76.260 135.980 76.460 ;
        RECT 131.240 76.120 132.760 76.260 ;
        RECT 133.080 76.120 135.980 76.260 ;
        RECT 107.230 75.920 107.550 75.980 ;
        RECT 108.625 75.920 108.915 75.965 ;
        RECT 107.230 75.780 108.915 75.920 ;
        RECT 107.230 75.720 107.550 75.780 ;
        RECT 108.625 75.735 108.915 75.780 ;
        RECT 119.665 75.920 119.955 75.965 ;
        RECT 121.490 75.920 121.810 75.980 ;
        RECT 119.665 75.780 121.810 75.920 ;
        RECT 119.665 75.735 119.955 75.780 ;
        RECT 121.490 75.720 121.810 75.780 ;
        RECT 127.010 75.920 127.330 75.980 ;
        RECT 131.625 75.920 131.915 75.965 ;
        RECT 127.010 75.780 131.915 75.920 ;
        RECT 132.620 75.920 132.760 76.120 ;
        RECT 141.360 75.980 141.500 76.460 ;
        RECT 142.205 76.460 143.430 76.600 ;
        RECT 142.205 76.415 142.495 76.460 ;
        RECT 143.110 76.400 143.430 76.460 ;
        RECT 143.585 76.415 143.875 76.645 ;
        RECT 143.660 76.260 143.800 76.415 ;
        RECT 142.740 76.120 143.800 76.260 ;
        RECT 142.740 75.980 142.880 76.120 ;
        RECT 134.845 75.920 135.135 75.965 ;
        RECT 132.620 75.780 135.135 75.920 ;
        RECT 127.010 75.720 127.330 75.780 ;
        RECT 131.625 75.735 131.915 75.780 ;
        RECT 134.845 75.735 135.135 75.780 ;
        RECT 137.145 75.920 137.435 75.965 ;
        RECT 138.970 75.920 139.290 75.980 ;
        RECT 137.145 75.780 139.290 75.920 ;
        RECT 137.145 75.735 137.435 75.780 ;
        RECT 138.970 75.720 139.290 75.780 ;
        RECT 141.270 75.720 141.590 75.980 ;
        RECT 141.730 75.720 142.050 75.980 ;
        RECT 142.650 75.720 142.970 75.980 ;
        RECT 145.410 75.720 145.730 75.980 ;
        RECT 146.790 75.720 147.110 75.980 ;
        RECT 152.900 75.580 153.380 80.540 ;
        RECT 91.060 75.100 153.380 75.580 ;
        RECT 105.850 74.900 106.170 74.960 ;
        RECT 115.510 74.900 115.830 74.960 ;
        RECT 105.850 74.760 115.830 74.900 ;
        RECT 105.850 74.700 106.170 74.760 ;
        RECT 115.510 74.700 115.830 74.760 ;
        RECT 118.730 74.900 119.050 74.960 ;
        RECT 119.665 74.900 119.955 74.945 ;
        RECT 118.730 74.760 119.955 74.900 ;
        RECT 118.730 74.700 119.050 74.760 ;
        RECT 119.665 74.715 119.955 74.760 ;
        RECT 130.690 74.700 131.010 74.960 ;
        RECT 138.970 74.700 139.290 74.960 ;
        RECT 141.270 74.700 141.590 74.960 ;
        RECT 146.790 74.700 147.110 74.960 ;
        RECT 105.355 74.560 105.645 74.605 ;
        RECT 107.245 74.560 107.535 74.605 ;
        RECT 110.365 74.560 110.655 74.605 ;
        RECT 105.355 74.420 110.655 74.560 ;
        RECT 105.355 74.375 105.645 74.420 ;
        RECT 107.245 74.375 107.535 74.420 ;
        RECT 110.365 74.375 110.655 74.420 ;
        RECT 119.190 74.560 119.510 74.620 ;
        RECT 126.105 74.560 126.395 74.605 ;
        RECT 135.750 74.560 136.070 74.620 ;
        RECT 139.060 74.560 139.200 74.700 ;
        RECT 142.650 74.560 142.970 74.620 ;
        RECT 119.190 74.420 126.395 74.560 ;
        RECT 119.190 74.360 119.510 74.420 ;
        RECT 126.105 74.375 126.395 74.420 ;
        RECT 132.160 74.420 139.200 74.560 ;
        RECT 141.820 74.420 142.970 74.560 ;
        RECT 104.485 74.220 104.775 74.265 ;
        RECT 116.445 74.220 116.735 74.265 ;
        RECT 118.270 74.220 118.590 74.280 ;
        RECT 104.485 74.080 111.140 74.220 ;
        RECT 104.485 74.035 104.775 74.080 ;
        RECT 111.000 73.940 111.140 74.080 ;
        RECT 116.445 74.080 118.590 74.220 ;
        RECT 116.445 74.035 116.735 74.080 ;
        RECT 118.270 74.020 118.590 74.080 ;
        RECT 121.045 74.220 121.335 74.265 ;
        RECT 132.160 74.220 132.300 74.420 ;
        RECT 135.750 74.360 136.070 74.420 ;
        RECT 138.050 74.220 138.370 74.280 ;
        RECT 121.045 74.080 122.640 74.220 ;
        RECT 121.045 74.035 121.335 74.080 ;
        RECT 122.500 73.940 122.640 74.080 ;
        RECT 131.700 74.080 132.300 74.220 ;
        RECT 133.770 74.080 138.370 74.220 ;
        RECT 104.950 73.880 105.240 73.925 ;
        RECT 106.785 73.880 107.075 73.925 ;
        RECT 110.365 73.880 110.655 73.925 ;
        RECT 104.950 73.740 110.655 73.880 ;
        RECT 104.950 73.695 105.240 73.740 ;
        RECT 106.785 73.695 107.075 73.740 ;
        RECT 110.365 73.695 110.655 73.740 ;
        RECT 110.910 73.680 111.230 73.940 ;
        RECT 105.865 73.540 106.155 73.585 ;
        RECT 107.230 73.540 107.550 73.600 ;
        RECT 105.865 73.400 107.550 73.540 ;
        RECT 105.865 73.355 106.155 73.400 ;
        RECT 107.230 73.340 107.550 73.400 ;
        RECT 108.145 73.540 108.795 73.585 ;
        RECT 109.070 73.540 109.390 73.600 ;
        RECT 111.445 73.585 111.735 73.900 ;
        RECT 115.985 73.695 116.275 73.925 ;
        RECT 111.445 73.540 112.035 73.585 ;
        RECT 108.145 73.400 112.035 73.540 ;
        RECT 108.145 73.355 108.795 73.400 ;
        RECT 109.070 73.340 109.390 73.400 ;
        RECT 111.745 73.355 112.035 73.400 ;
        RECT 114.605 73.540 114.895 73.585 ;
        RECT 116.060 73.540 116.200 73.695 ;
        RECT 120.570 73.680 120.890 73.940 ;
        RECT 121.490 73.680 121.810 73.940 ;
        RECT 121.950 73.680 122.270 73.940 ;
        RECT 122.410 73.680 122.730 73.940 ;
        RECT 131.700 73.925 131.840 74.080 ;
        RECT 133.770 73.975 133.910 74.080 ;
        RECT 138.050 74.020 138.370 74.080 ;
        RECT 122.960 73.740 131.380 73.880 ;
        RECT 121.580 73.540 121.720 73.680 ;
        RECT 122.960 73.540 123.100 73.740 ;
        RECT 114.605 73.400 123.100 73.540 ;
        RECT 114.605 73.355 114.895 73.400 ;
        RECT 127.010 73.340 127.330 73.600 ;
        RECT 127.470 73.540 127.790 73.600 ;
        RECT 127.945 73.540 128.235 73.585 ;
        RECT 127.470 73.400 128.235 73.540 ;
        RECT 131.240 73.540 131.380 73.740 ;
        RECT 131.625 73.695 131.915 73.925 ;
        RECT 132.085 73.695 132.375 73.925 ;
        RECT 133.005 73.695 133.295 73.925 ;
        RECT 133.515 73.790 133.910 73.975 ;
        RECT 133.515 73.745 133.805 73.790 ;
        RECT 132.160 73.540 132.300 73.695 ;
        RECT 131.240 73.400 132.300 73.540 ;
        RECT 133.080 73.540 133.220 73.695 ;
        RECT 137.590 73.680 137.910 73.940 ;
        RECT 141.270 73.880 141.590 73.940 ;
        RECT 141.820 73.925 141.960 74.420 ;
        RECT 142.650 74.360 142.970 74.420 ;
        RECT 146.880 74.220 147.020 74.700 ;
        RECT 142.280 74.080 144.720 74.220 ;
        RECT 142.280 73.940 142.420 74.080 ;
        RECT 141.745 73.880 142.035 73.925 ;
        RECT 141.270 73.740 142.035 73.880 ;
        RECT 141.270 73.680 141.590 73.740 ;
        RECT 141.745 73.695 142.035 73.740 ;
        RECT 142.190 73.680 142.510 73.940 ;
        RECT 142.665 73.880 142.955 73.925 ;
        RECT 143.110 73.880 143.430 73.940 ;
        RECT 142.665 73.740 143.430 73.880 ;
        RECT 142.665 73.695 142.955 73.740 ;
        RECT 143.110 73.680 143.430 73.740 ;
        RECT 143.570 73.680 143.890 73.940 ;
        RECT 133.450 73.540 133.770 73.600 ;
        RECT 133.080 73.400 133.770 73.540 ;
        RECT 127.470 73.340 127.790 73.400 ;
        RECT 127.945 73.355 128.235 73.400 ;
        RECT 117.825 73.200 118.115 73.245 ;
        RECT 118.730 73.200 119.050 73.260 ;
        RECT 117.825 73.060 119.050 73.200 ;
        RECT 132.160 73.200 132.300 73.400 ;
        RECT 133.450 73.340 133.770 73.400 ;
        RECT 135.290 73.200 135.610 73.260 ;
        RECT 137.680 73.200 137.820 73.680 ;
        RECT 144.045 73.540 144.335 73.585 ;
        RECT 140.900 73.400 144.335 73.540 ;
        RECT 144.580 73.540 144.720 74.080 ;
        RECT 145.500 74.080 147.020 74.220 ;
        RECT 145.500 73.925 145.640 74.080 ;
        RECT 145.425 73.695 145.715 73.925 ;
        RECT 145.870 73.680 146.190 73.940 ;
        RECT 146.330 73.680 146.650 73.940 ;
        RECT 147.265 73.695 147.555 73.925 ;
        RECT 145.960 73.540 146.100 73.680 ;
        RECT 144.580 73.400 146.100 73.540 ;
        RECT 140.900 73.260 141.040 73.400 ;
        RECT 144.045 73.355 144.335 73.400 ;
        RECT 132.160 73.060 137.820 73.200 ;
        RECT 117.825 73.015 118.115 73.060 ;
        RECT 118.730 73.000 119.050 73.060 ;
        RECT 135.290 73.000 135.610 73.060 ;
        RECT 140.810 73.000 141.130 73.260 ;
        RECT 143.110 73.000 143.430 73.260 ;
        RECT 145.870 73.200 146.190 73.260 ;
        RECT 147.340 73.200 147.480 73.695 ;
        RECT 145.870 73.060 147.480 73.200 ;
        RECT 145.870 73.000 146.190 73.060 ;
        RECT 88.980 72.380 152.240 72.860 ;
        RECT 88.980 67.420 89.460 72.380 ;
        RECT 109.070 71.980 109.390 72.240 ;
        RECT 115.050 72.180 115.370 72.240 ;
        RECT 117.365 72.180 117.655 72.225 ;
        RECT 125.645 72.180 125.935 72.225 ;
        RECT 136.670 72.180 136.990 72.240 ;
        RECT 115.050 72.040 117.655 72.180 ;
        RECT 115.050 71.980 115.370 72.040 ;
        RECT 117.365 71.995 117.655 72.040 ;
        RECT 118.360 72.040 125.935 72.180 ;
        RECT 118.360 71.840 118.500 72.040 ;
        RECT 125.645 71.995 125.935 72.040 ;
        RECT 134.000 72.040 136.990 72.180 ;
        RECT 115.140 71.700 118.500 71.840 ;
        RECT 118.730 71.840 119.050 71.900 ;
        RECT 119.665 71.840 119.955 71.885 ;
        RECT 127.470 71.840 127.790 71.900 ;
        RECT 133.465 71.840 133.755 71.885 ;
        RECT 118.730 71.700 119.955 71.840 ;
        RECT 108.625 71.500 108.915 71.545 ;
        RECT 109.530 71.500 109.850 71.560 ;
        RECT 112.750 71.500 113.070 71.560 ;
        RECT 115.140 71.545 115.280 71.700 ;
        RECT 118.730 71.640 119.050 71.700 ;
        RECT 119.665 71.655 119.955 71.700 ;
        RECT 120.660 71.700 126.320 71.840 ;
        RECT 120.660 71.560 120.800 71.700 ;
        RECT 108.625 71.360 113.070 71.500 ;
        RECT 108.625 71.315 108.915 71.360 ;
        RECT 109.530 71.300 109.850 71.360 ;
        RECT 112.750 71.300 113.070 71.360 ;
        RECT 115.065 71.315 115.355 71.545 ;
        RECT 115.985 71.315 116.275 71.545 ;
        RECT 116.445 71.500 116.735 71.545 ;
        RECT 116.445 71.360 118.500 71.500 ;
        RECT 116.445 71.315 116.735 71.360 ;
        RECT 115.050 70.280 115.370 70.540 ;
        RECT 116.060 70.480 116.200 71.315 ;
        RECT 118.360 71.220 118.500 71.360 ;
        RECT 120.570 71.300 120.890 71.560 ;
        RECT 126.180 71.545 126.320 71.700 ;
        RECT 127.470 71.700 133.755 71.840 ;
        RECT 127.470 71.640 127.790 71.700 ;
        RECT 133.465 71.655 133.755 71.700 ;
        RECT 124.725 71.500 125.015 71.545 ;
        RECT 125.185 71.500 125.475 71.545 ;
        RECT 124.725 71.360 125.475 71.500 ;
        RECT 124.725 71.315 125.015 71.360 ;
        RECT 125.185 71.315 125.475 71.360 ;
        RECT 126.105 71.315 126.395 71.545 ;
        RECT 126.565 71.500 126.855 71.545 ;
        RECT 127.010 71.500 127.330 71.560 ;
        RECT 126.565 71.360 127.330 71.500 ;
        RECT 126.565 71.315 126.855 71.360 ;
        RECT 127.010 71.300 127.330 71.360 ;
        RECT 127.945 71.500 128.235 71.545 ;
        RECT 134.000 71.500 134.140 72.040 ;
        RECT 136.670 71.980 136.990 72.040 ;
        RECT 138.970 71.980 139.290 72.240 ;
        RECT 140.350 72.180 140.670 72.240 ;
        RECT 144.965 72.180 145.255 72.225 ;
        RECT 145.410 72.180 145.730 72.240 ;
        RECT 140.350 72.040 143.800 72.180 ;
        RECT 140.350 71.980 140.670 72.040 ;
        RECT 143.660 71.840 143.800 72.040 ;
        RECT 144.965 72.040 145.730 72.180 ;
        RECT 144.965 71.995 145.255 72.040 ;
        RECT 145.410 71.980 145.730 72.040 ;
        RECT 148.630 71.840 148.950 71.900 ;
        RECT 135.380 71.700 143.340 71.840 ;
        RECT 143.660 71.700 148.950 71.840 ;
        RECT 127.945 71.360 134.140 71.500 ;
        RECT 127.945 71.315 128.235 71.360 ;
        RECT 134.370 71.300 134.690 71.560 ;
        RECT 135.380 71.545 135.520 71.700 ;
        RECT 143.200 71.560 143.340 71.700 ;
        RECT 148.630 71.640 148.950 71.700 ;
        RECT 135.305 71.315 135.595 71.545 ;
        RECT 135.765 71.315 136.055 71.545 ;
        RECT 118.270 70.960 118.590 71.220 ;
        RECT 121.965 71.160 122.255 71.205 ;
        RECT 122.410 71.160 122.730 71.220 ;
        RECT 135.840 71.160 135.980 71.315 ;
        RECT 137.590 71.300 137.910 71.560 ;
        RECT 139.445 71.500 139.735 71.545 ;
        RECT 139.445 71.360 141.500 71.500 ;
        RECT 139.445 71.315 139.735 71.360 ;
        RECT 139.905 71.160 140.195 71.205 ;
        RECT 140.350 71.160 140.670 71.220 ;
        RECT 121.965 71.020 122.730 71.160 ;
        RECT 121.965 70.975 122.255 71.020 ;
        RECT 122.410 70.960 122.730 71.020 ;
        RECT 126.180 71.020 139.660 71.160 ;
        RECT 117.825 70.820 118.115 70.865 ;
        RECT 119.190 70.820 119.510 70.880 ;
        RECT 117.825 70.680 119.510 70.820 ;
        RECT 117.825 70.635 118.115 70.680 ;
        RECT 119.190 70.620 119.510 70.680 ;
        RECT 126.180 70.480 126.320 71.020 ;
        RECT 134.845 70.820 135.135 70.865 ;
        RECT 138.510 70.820 138.830 70.880 ;
        RECT 134.845 70.680 138.830 70.820 ;
        RECT 139.520 70.820 139.660 71.020 ;
        RECT 139.905 71.020 140.670 71.160 ;
        RECT 139.905 70.975 140.195 71.020 ;
        RECT 140.350 70.960 140.670 71.020 ;
        RECT 140.810 70.820 141.130 70.880 ;
        RECT 141.360 70.865 141.500 71.360 ;
        RECT 143.110 71.300 143.430 71.560 ;
        RECT 145.870 71.500 146.190 71.560 ;
        RECT 146.790 71.500 147.110 71.560 ;
        RECT 145.870 71.360 147.110 71.500 ;
        RECT 145.870 71.300 146.190 71.360 ;
        RECT 146.790 71.300 147.110 71.360 ;
        RECT 147.250 71.500 147.570 71.560 ;
        RECT 149.105 71.500 149.395 71.545 ;
        RECT 147.250 71.360 149.395 71.500 ;
        RECT 147.250 71.300 147.570 71.360 ;
        RECT 149.105 71.315 149.395 71.360 ;
        RECT 142.650 71.160 142.970 71.220 ;
        RECT 143.570 71.160 143.890 71.220 ;
        RECT 142.650 71.020 146.100 71.160 ;
        RECT 142.650 70.960 142.970 71.020 ;
        RECT 143.570 70.960 143.890 71.020 ;
        RECT 139.520 70.680 141.130 70.820 ;
        RECT 134.845 70.635 135.135 70.680 ;
        RECT 138.510 70.620 138.830 70.680 ;
        RECT 140.810 70.620 141.130 70.680 ;
        RECT 141.285 70.635 141.575 70.865 ;
        RECT 142.205 70.820 142.495 70.865 ;
        RECT 143.110 70.820 143.430 70.880 ;
        RECT 145.960 70.865 146.100 71.020 ;
        RECT 150.470 70.960 150.790 71.220 ;
        RECT 142.205 70.680 143.430 70.820 ;
        RECT 142.205 70.635 142.495 70.680 ;
        RECT 116.060 70.340 126.320 70.480 ;
        RECT 126.565 70.480 126.855 70.525 ;
        RECT 127.470 70.480 127.790 70.540 ;
        RECT 126.565 70.340 127.790 70.480 ;
        RECT 126.565 70.295 126.855 70.340 ;
        RECT 127.470 70.280 127.790 70.340 ;
        RECT 133.450 70.480 133.770 70.540 ;
        RECT 137.145 70.480 137.435 70.525 ;
        RECT 133.450 70.340 137.435 70.480 ;
        RECT 133.450 70.280 133.770 70.340 ;
        RECT 137.145 70.295 137.435 70.340 ;
        RECT 140.350 70.480 140.670 70.540 ;
        RECT 141.360 70.480 141.500 70.635 ;
        RECT 143.110 70.620 143.430 70.680 ;
        RECT 145.885 70.635 146.175 70.865 ;
        RECT 140.350 70.340 141.500 70.480 ;
        RECT 144.965 70.480 145.255 70.525 ;
        RECT 145.410 70.480 145.730 70.540 ;
        RECT 144.965 70.340 145.730 70.480 ;
        RECT 140.350 70.280 140.670 70.340 ;
        RECT 144.965 70.295 145.255 70.340 ;
        RECT 145.410 70.280 145.730 70.340 ;
        RECT 152.900 70.140 153.380 75.100 ;
        RECT 91.060 69.660 153.380 70.140 ;
        RECT 118.270 69.460 118.590 69.520 ;
        RECT 120.585 69.460 120.875 69.505 ;
        RECT 118.270 69.320 120.875 69.460 ;
        RECT 118.270 69.260 118.590 69.320 ;
        RECT 120.585 69.275 120.875 69.320 ;
        RECT 134.370 69.260 134.690 69.520 ;
        RECT 135.290 69.260 135.610 69.520 ;
        RECT 138.050 69.260 138.370 69.520 ;
        RECT 138.510 69.460 138.830 69.520 ;
        RECT 139.905 69.460 140.195 69.505 ;
        RECT 138.510 69.320 140.195 69.460 ;
        RECT 138.510 69.260 138.830 69.320 ;
        RECT 139.905 69.275 140.195 69.320 ;
        RECT 140.350 69.460 140.670 69.520 ;
        RECT 144.030 69.460 144.350 69.520 ;
        RECT 140.350 69.320 144.350 69.460 ;
        RECT 140.350 69.260 140.670 69.320 ;
        RECT 144.030 69.260 144.350 69.320 ;
        RECT 145.885 69.460 146.175 69.505 ;
        RECT 146.330 69.460 146.650 69.520 ;
        RECT 145.885 69.320 146.650 69.460 ;
        RECT 145.885 69.275 146.175 69.320 ;
        RECT 146.330 69.260 146.650 69.320 ;
        RECT 147.265 69.275 147.555 69.505 ;
        RECT 111.795 69.120 112.085 69.165 ;
        RECT 113.685 69.120 113.975 69.165 ;
        RECT 116.805 69.120 117.095 69.165 ;
        RECT 111.795 68.980 117.095 69.120 ;
        RECT 111.795 68.935 112.085 68.980 ;
        RECT 113.685 68.935 113.975 68.980 ;
        RECT 116.805 68.935 117.095 68.980 ;
        RECT 133.925 69.120 134.215 69.165 ;
        RECT 135.380 69.120 135.520 69.260 ;
        RECT 133.925 68.980 135.520 69.120 ;
        RECT 133.925 68.935 134.215 68.980 ;
        RECT 137.590 68.920 137.910 69.180 ;
        RECT 110.910 68.580 111.230 68.840 ;
        RECT 112.305 68.780 112.595 68.825 ;
        RECT 115.050 68.780 115.370 68.840 ;
        RECT 112.305 68.640 115.370 68.780 ;
        RECT 112.305 68.595 112.595 68.640 ;
        RECT 115.050 68.580 115.370 68.640 ;
        RECT 119.665 68.780 119.955 68.825 ;
        RECT 132.085 68.780 132.375 68.825 ;
        RECT 137.680 68.780 137.820 68.920 ;
        RECT 140.810 68.780 141.130 68.840 ;
        RECT 119.665 68.640 122.640 68.780 ;
        RECT 119.665 68.595 119.955 68.640 ;
        RECT 122.500 68.500 122.640 68.640 ;
        RECT 132.085 68.640 141.130 68.780 ;
        RECT 132.085 68.595 132.375 68.640 ;
        RECT 102.185 68.440 102.475 68.485 ;
        RECT 103.550 68.440 103.870 68.500 ;
        RECT 102.185 68.300 103.870 68.440 ;
        RECT 102.185 68.255 102.475 68.300 ;
        RECT 103.550 68.240 103.870 68.300 ;
        RECT 111.390 68.440 111.680 68.485 ;
        RECT 113.225 68.440 113.515 68.485 ;
        RECT 116.805 68.440 117.095 68.485 ;
        RECT 111.390 68.300 117.095 68.440 ;
        RECT 111.390 68.255 111.680 68.300 ;
        RECT 113.225 68.255 113.515 68.300 ;
        RECT 116.805 68.255 117.095 68.300 ;
        RECT 115.050 68.145 115.370 68.160 ;
        RECT 114.585 68.100 115.370 68.145 ;
        RECT 117.885 68.145 118.175 68.460 ;
        RECT 121.505 68.440 121.795 68.485 ;
        RECT 121.120 68.300 121.795 68.440 ;
        RECT 117.885 68.100 118.475 68.145 ;
        RECT 114.585 67.960 118.475 68.100 ;
        RECT 114.585 67.915 115.370 67.960 ;
        RECT 118.185 67.915 118.475 67.960 ;
        RECT 115.050 67.900 115.370 67.915 ;
        RECT 121.120 67.820 121.260 68.300 ;
        RECT 121.505 68.255 121.795 68.300 ;
        RECT 122.410 68.240 122.730 68.500 ;
        RECT 134.920 68.485 135.060 68.640 ;
        RECT 140.810 68.580 141.130 68.640 ;
        RECT 143.570 68.580 143.890 68.840 ;
        RECT 145.410 68.780 145.730 68.840 ;
        RECT 146.345 68.780 146.635 68.825 ;
        RECT 145.410 68.640 146.635 68.780 ;
        RECT 145.410 68.580 145.730 68.640 ;
        RECT 146.345 68.595 146.635 68.640 ;
        RECT 134.845 68.255 135.135 68.485 ;
        RECT 137.605 68.440 137.895 68.485 ;
        RECT 137.220 68.300 137.895 68.440 ;
        RECT 100.330 67.760 100.650 67.820 ;
        RECT 101.265 67.760 101.555 67.805 ;
        RECT 100.330 67.620 101.555 67.760 ;
        RECT 100.330 67.560 100.650 67.620 ;
        RECT 101.265 67.575 101.555 67.620 ;
        RECT 121.030 67.560 121.350 67.820 ;
        RECT 135.290 67.760 135.610 67.820 ;
        RECT 137.220 67.805 137.360 68.300 ;
        RECT 137.605 68.255 137.895 68.300 ;
        RECT 141.730 68.440 142.050 68.500 ;
        RECT 142.665 68.440 142.955 68.485 ;
        RECT 141.730 68.300 142.955 68.440 ;
        RECT 141.730 68.240 142.050 68.300 ;
        RECT 142.665 68.255 142.955 68.300 ;
        RECT 143.110 68.240 143.430 68.500 ;
        RECT 143.660 68.440 143.800 68.580 ;
        RECT 144.990 68.450 145.280 68.485 ;
        RECT 144.580 68.440 145.280 68.450 ;
        RECT 143.660 68.310 145.280 68.440 ;
        RECT 143.660 68.300 144.720 68.310 ;
        RECT 144.990 68.255 145.280 68.310 ;
        RECT 144.045 67.915 144.335 68.145 ;
        RECT 144.505 67.915 144.795 68.145 ;
        RECT 147.340 68.100 147.480 69.275 ;
        RECT 148.630 68.240 148.950 68.500 ;
        RECT 145.500 67.960 147.480 68.100 ;
        RECT 137.145 67.760 137.435 67.805 ;
        RECT 135.290 67.620 137.435 67.760 ;
        RECT 135.290 67.560 135.610 67.620 ;
        RECT 137.145 67.575 137.435 67.620 ;
        RECT 142.650 67.760 142.970 67.820 ;
        RECT 144.120 67.760 144.260 67.915 ;
        RECT 142.650 67.620 144.260 67.760 ;
        RECT 144.580 67.760 144.720 67.915 ;
        RECT 145.500 67.820 145.640 67.960 ;
        RECT 144.950 67.760 145.270 67.820 ;
        RECT 144.580 67.620 145.270 67.760 ;
        RECT 142.650 67.560 142.970 67.620 ;
        RECT 144.950 67.560 145.270 67.620 ;
        RECT 145.410 67.560 145.730 67.820 ;
        RECT 145.870 67.760 146.190 67.820 ;
        RECT 147.250 67.760 147.570 67.820 ;
        RECT 145.870 67.620 147.570 67.760 ;
        RECT 145.870 67.560 146.190 67.620 ;
        RECT 147.250 67.560 147.570 67.620 ;
        RECT 88.980 66.940 152.240 67.420 ;
        RECT 31.665 66.710 34.250 66.735 ;
        RECT 31.665 66.660 32.005 66.710 ;
        RECT 33.840 66.655 34.250 66.710 ;
        RECT 21.870 65.390 22.100 66.390 ;
        RECT 22.310 65.390 22.540 66.390 ;
        RECT 23.510 65.350 23.740 66.350 ;
        RECT 23.950 65.350 24.180 66.350 ;
        RECT 24.390 65.350 24.620 66.350 ;
        RECT 25.040 65.350 25.270 66.350 ;
        RECT 25.480 65.350 25.710 66.350 ;
        RECT 25.920 65.350 26.150 66.350 ;
        RECT 26.530 65.350 26.760 66.350 ;
        RECT 26.970 65.350 27.200 66.350 ;
        RECT 28.840 65.350 29.070 66.350 ;
        RECT 29.280 65.350 29.510 66.350 ;
        RECT 29.720 65.350 29.950 66.350 ;
        RECT 30.370 65.350 30.600 66.350 ;
        RECT 30.810 65.350 31.040 66.350 ;
        RECT 31.250 65.350 31.480 66.350 ;
        RECT 32.065 65.290 32.295 66.290 ;
        RECT 32.505 65.290 32.735 66.290 ;
        RECT 33.115 65.290 33.345 66.290 ;
        RECT 33.555 65.290 33.785 66.290 ;
        RECT 35.135 65.595 35.590 65.975 ;
        RECT 21.870 63.720 22.100 64.720 ;
        RECT 22.310 63.720 22.540 64.720 ;
        RECT 18.930 63.285 19.550 63.720 ;
        RECT 23.510 63.400 23.740 64.400 ;
        RECT 23.950 63.400 24.180 64.400 ;
        RECT 24.390 63.400 24.620 64.400 ;
        RECT 25.040 63.400 25.270 64.400 ;
        RECT 25.480 63.400 25.710 64.400 ;
        RECT 25.920 63.400 26.150 64.400 ;
        RECT 26.530 63.680 26.760 64.680 ;
        RECT 26.970 63.680 27.200 64.680 ;
        RECT 21.415 61.730 21.845 62.240 ;
        RECT 6.080 56.695 6.330 58.800 ;
        RECT 21.440 58.500 21.795 61.730 ;
        RECT 8.125 58.175 21.800 58.500 ;
        RECT 7.365 57.690 21.800 58.175 ;
        RECT 7.365 57.315 8.285 57.690 ;
        RECT 22.730 56.360 23.980 57.440 ;
        RECT 6.080 53.540 6.330 55.645 ;
        RECT 6.020 51.220 6.380 51.390 ;
        RECT 24.420 51.220 24.590 63.400 ;
        RECT 27.550 63.225 28.240 63.780 ;
        RECT 28.840 63.400 29.070 64.400 ;
        RECT 29.280 63.400 29.510 64.400 ;
        RECT 29.720 63.400 29.950 64.400 ;
        RECT 30.370 63.400 30.600 64.400 ;
        RECT 30.810 63.400 31.040 64.400 ;
        RECT 31.250 63.400 31.480 64.400 ;
        RECT 32.065 63.620 32.295 64.620 ;
        RECT 32.505 63.620 32.735 64.620 ;
        RECT 33.115 63.620 33.345 64.620 ;
        RECT 33.555 63.620 33.785 64.620 ;
        RECT 34.430 64.585 34.980 65.080 ;
        RECT 34.455 64.580 34.835 64.585 ;
        RECT 31.040 62.610 31.455 62.650 ;
        RECT 31.040 62.450 56.015 62.610 ;
        RECT 31.040 62.385 31.455 62.450 ;
        RECT 32.650 61.770 32.930 61.850 ;
        RECT 53.130 61.770 54.030 61.775 ;
        RECT 32.650 61.600 54.030 61.770 ;
        RECT 32.650 61.535 32.930 61.600 ;
        RECT 53.130 61.090 54.030 61.600 ;
        RECT 24.890 59.335 25.425 59.755 ;
        RECT 6.020 51.050 24.590 51.220 ;
        RECT 25.005 51.165 25.285 59.335 ;
        RECT 28.685 59.095 29.310 59.605 ;
        RECT 29.750 59.505 30.145 59.570 ;
        RECT 33.990 59.505 34.890 59.725 ;
        RECT 29.750 59.265 34.890 59.505 ;
        RECT 29.750 59.205 30.145 59.265 ;
        RECT 28.690 59.090 29.305 59.095 ;
        RECT 33.990 59.080 34.890 59.265 ;
        RECT 26.380 57.705 27.105 58.735 ;
        RECT 55.855 57.505 56.015 62.450 ;
        RECT 88.980 61.980 89.460 66.940 ;
        RECT 109.530 66.740 109.850 66.800 ;
        RECT 115.050 66.740 115.370 66.800 ;
        RECT 122.410 66.740 122.730 66.800 ;
        RECT 138.050 66.740 138.370 66.800 ;
        RECT 109.530 66.600 114.820 66.740 ;
        RECT 109.530 66.540 109.850 66.600 ;
        RECT 99.885 66.400 100.175 66.445 ;
        RECT 100.330 66.400 100.650 66.460 ;
        RECT 99.885 66.260 100.650 66.400 ;
        RECT 99.885 66.215 100.175 66.260 ;
        RECT 100.330 66.200 100.650 66.260 ;
        RECT 102.165 66.400 102.815 66.445 ;
        RECT 105.765 66.400 106.055 66.445 ;
        RECT 108.625 66.400 108.915 66.445 ;
        RECT 102.165 66.260 108.915 66.400 ;
        RECT 102.165 66.215 102.815 66.260 ;
        RECT 105.465 66.215 106.055 66.260 ;
        RECT 108.625 66.215 108.915 66.260 ;
        RECT 98.970 66.060 99.260 66.105 ;
        RECT 100.805 66.060 101.095 66.105 ;
        RECT 104.385 66.060 104.675 66.105 ;
        RECT 98.970 65.920 104.675 66.060 ;
        RECT 98.970 65.875 99.260 65.920 ;
        RECT 100.805 65.875 101.095 65.920 ;
        RECT 104.385 65.875 104.675 65.920 ;
        RECT 105.465 65.900 105.755 66.215 ;
        RECT 109.085 66.060 109.375 66.105 ;
        RECT 106.860 65.920 109.375 66.060 ;
        RECT 114.680 66.060 114.820 66.600 ;
        RECT 115.050 66.600 115.740 66.740 ;
        RECT 115.050 66.540 115.370 66.600 ;
        RECT 115.600 66.445 115.740 66.600 ;
        RECT 122.410 66.600 138.370 66.740 ;
        RECT 122.410 66.540 122.730 66.600 ;
        RECT 127.930 66.445 128.250 66.460 ;
        RECT 115.525 66.215 115.815 66.445 ;
        RECT 127.925 66.400 128.575 66.445 ;
        RECT 131.525 66.400 131.815 66.445 ;
        RECT 127.925 66.260 131.815 66.400 ;
        RECT 127.925 66.215 128.575 66.260 ;
        RECT 131.225 66.215 131.815 66.260 ;
        RECT 127.930 66.200 128.250 66.215 ;
        RECT 115.065 66.060 115.355 66.105 ;
        RECT 114.680 65.920 115.355 66.060 ;
        RECT 98.505 65.535 98.795 65.765 ;
        RECT 98.580 65.040 98.720 65.535 ;
        RECT 99.375 65.380 99.665 65.425 ;
        RECT 101.265 65.380 101.555 65.425 ;
        RECT 104.385 65.380 104.675 65.425 ;
        RECT 99.375 65.240 104.675 65.380 ;
        RECT 99.375 65.195 99.665 65.240 ;
        RECT 101.265 65.195 101.555 65.240 ;
        RECT 104.385 65.195 104.675 65.240 ;
        RECT 101.710 65.040 102.030 65.100 ;
        RECT 98.580 64.900 102.030 65.040 ;
        RECT 101.710 64.840 102.030 64.900 ;
        RECT 103.090 65.040 103.410 65.100 ;
        RECT 106.860 65.040 107.000 65.920 ;
        RECT 109.085 65.875 109.375 65.920 ;
        RECT 115.065 65.875 115.355 65.920 ;
        RECT 122.885 65.875 123.175 66.105 ;
        RECT 109.160 65.720 109.300 65.875 ;
        RECT 122.960 65.720 123.100 65.875 ;
        RECT 124.250 65.860 124.570 66.120 ;
        RECT 124.730 66.060 125.020 66.105 ;
        RECT 126.565 66.060 126.855 66.105 ;
        RECT 130.145 66.060 130.435 66.105 ;
        RECT 124.730 65.920 130.435 66.060 ;
        RECT 124.730 65.875 125.020 65.920 ;
        RECT 126.565 65.875 126.855 65.920 ;
        RECT 130.145 65.875 130.435 65.920 ;
        RECT 131.225 65.900 131.515 66.215 ;
        RECT 134.000 66.105 134.140 66.600 ;
        RECT 138.050 66.540 138.370 66.600 ;
        RECT 143.110 66.540 143.430 66.800 ;
        RECT 135.305 66.400 135.595 66.445 ;
        RECT 143.200 66.400 143.340 66.540 ;
        RECT 135.305 66.260 143.340 66.400 ;
        RECT 135.305 66.215 135.595 66.260 ;
        RECT 133.925 65.875 134.215 66.105 ;
        RECT 134.370 65.860 134.690 66.120 ;
        RECT 139.445 66.060 139.735 66.105 ;
        RECT 139.890 66.060 140.210 66.120 ;
        RECT 134.920 65.920 140.210 66.060 ;
        RECT 109.160 65.580 123.100 65.720 ;
        RECT 125.645 65.720 125.935 65.765 ;
        RECT 127.470 65.720 127.790 65.780 ;
        RECT 125.645 65.580 127.790 65.720 ;
        RECT 125.645 65.535 125.935 65.580 ;
        RECT 127.470 65.520 127.790 65.580 ;
        RECT 133.005 65.720 133.295 65.765 ;
        RECT 134.920 65.720 135.060 65.920 ;
        RECT 139.445 65.875 139.735 65.920 ;
        RECT 139.890 65.860 140.210 65.920 ;
        RECT 141.745 66.060 142.035 66.105 ;
        RECT 144.030 66.060 144.350 66.120 ;
        RECT 144.505 66.060 144.795 66.105 ;
        RECT 145.410 66.060 145.730 66.120 ;
        RECT 141.745 65.920 145.730 66.060 ;
        RECT 141.745 65.875 142.035 65.920 ;
        RECT 144.030 65.860 144.350 65.920 ;
        RECT 144.505 65.875 144.795 65.920 ;
        RECT 145.410 65.860 145.730 65.920 ;
        RECT 145.870 65.860 146.190 66.120 ;
        RECT 133.005 65.580 135.060 65.720 ;
        RECT 133.005 65.535 133.295 65.580 ;
        RECT 135.290 65.520 135.610 65.780 ;
        RECT 140.365 65.720 140.655 65.765 ;
        RECT 142.190 65.720 142.510 65.780 ;
        RECT 144.965 65.720 145.255 65.765 ;
        RECT 140.365 65.580 145.255 65.720 ;
        RECT 140.365 65.535 140.655 65.580 ;
        RECT 142.190 65.520 142.510 65.580 ;
        RECT 144.965 65.535 145.255 65.580 ;
        RECT 125.135 65.380 125.425 65.425 ;
        RECT 127.025 65.380 127.315 65.425 ;
        RECT 130.145 65.380 130.435 65.425 ;
        RECT 125.135 65.240 130.435 65.380 ;
        RECT 125.135 65.195 125.425 65.240 ;
        RECT 127.025 65.195 127.315 65.240 ;
        RECT 130.145 65.195 130.435 65.240 ;
        RECT 139.905 65.380 140.195 65.425 ;
        RECT 141.270 65.380 141.590 65.440 ;
        RECT 145.960 65.380 146.100 65.860 ;
        RECT 139.905 65.240 146.100 65.380 ;
        RECT 139.905 65.195 140.195 65.240 ;
        RECT 141.270 65.180 141.590 65.240 ;
        RECT 103.090 64.900 107.000 65.040 ;
        RECT 103.090 64.840 103.410 64.900 ;
        RECT 107.230 64.840 107.550 65.100 ;
        RECT 122.410 64.840 122.730 65.100 ;
        RECT 138.050 64.840 138.370 65.100 ;
        RECT 140.810 65.040 141.130 65.100 ;
        RECT 142.650 65.040 142.970 65.100 ;
        RECT 140.810 64.900 142.970 65.040 ;
        RECT 140.810 64.840 141.130 64.900 ;
        RECT 142.650 64.840 142.970 64.900 ;
        RECT 143.110 65.040 143.430 65.100 ;
        RECT 143.585 65.040 143.875 65.085 ;
        RECT 143.110 64.900 143.875 65.040 ;
        RECT 143.110 64.840 143.430 64.900 ;
        RECT 143.585 64.855 143.875 64.900 ;
        RECT 144.030 65.040 144.350 65.100 ;
        RECT 145.885 65.040 146.175 65.085 ;
        RECT 150.930 65.040 151.250 65.100 ;
        RECT 144.030 64.900 151.250 65.040 ;
        RECT 144.030 64.840 144.350 64.900 ;
        RECT 145.885 64.855 146.175 64.900 ;
        RECT 150.930 64.840 151.250 64.900 ;
        RECT 152.900 64.700 153.380 69.660 ;
        RECT 91.060 64.220 153.380 64.700 ;
        RECT 101.710 64.020 102.030 64.080 ;
        RECT 110.910 64.020 111.230 64.080 ;
        RECT 101.710 63.880 111.230 64.020 ;
        RECT 101.710 63.820 102.030 63.880 ;
        RECT 110.910 63.820 111.230 63.880 ;
        RECT 122.410 63.820 122.730 64.080 ;
        RECT 127.025 64.020 127.315 64.065 ;
        RECT 127.930 64.020 128.250 64.080 ;
        RECT 127.025 63.880 128.250 64.020 ;
        RECT 127.025 63.835 127.315 63.880 ;
        RECT 127.930 63.820 128.250 63.880 ;
        RECT 146.330 64.020 146.650 64.080 ;
        RECT 146.805 64.020 147.095 64.065 ;
        RECT 146.330 63.880 147.095 64.020 ;
        RECT 146.330 63.820 146.650 63.880 ;
        RECT 146.805 63.835 147.095 63.880 ;
        RECT 95.845 63.680 96.135 63.725 ;
        RECT 98.965 63.680 99.255 63.725 ;
        RECT 100.855 63.680 101.145 63.725 ;
        RECT 95.845 63.540 101.145 63.680 ;
        RECT 95.845 63.495 96.135 63.540 ;
        RECT 98.965 63.495 99.255 63.540 ;
        RECT 100.855 63.495 101.145 63.540 ;
        RECT 101.800 63.385 101.940 63.820 ;
        RECT 110.465 63.680 110.755 63.725 ;
        RECT 113.635 63.680 113.925 63.725 ;
        RECT 115.525 63.680 115.815 63.725 ;
        RECT 118.645 63.680 118.935 63.725 ;
        RECT 122.500 63.680 122.640 63.820 ;
        RECT 143.110 63.680 143.430 63.740 ;
        RECT 107.780 63.540 112.520 63.680 ;
        RECT 101.725 63.155 102.015 63.385 ;
        RECT 106.660 63.340 106.950 63.385 ;
        RECT 107.230 63.340 107.550 63.400 ;
        RECT 106.660 63.200 107.550 63.340 ;
        RECT 106.660 63.155 106.950 63.200 ;
        RECT 107.230 63.140 107.550 63.200 ;
        RECT 107.780 63.045 107.920 63.540 ;
        RECT 110.465 63.495 110.755 63.540 ;
        RECT 94.765 62.705 95.055 63.020 ;
        RECT 95.845 63.000 96.135 63.045 ;
        RECT 99.425 63.000 99.715 63.045 ;
        RECT 101.260 63.000 101.550 63.045 ;
        RECT 95.845 62.860 101.550 63.000 ;
        RECT 95.845 62.815 96.135 62.860 ;
        RECT 99.425 62.815 99.715 62.860 ;
        RECT 101.260 62.815 101.550 62.860 ;
        RECT 103.105 62.815 103.395 63.045 ;
        RECT 107.705 62.815 107.995 63.045 ;
        RECT 109.085 63.000 109.375 63.045 ;
        RECT 109.085 62.860 112.060 63.000 ;
        RECT 109.085 62.815 109.375 62.860 ;
        RECT 94.465 62.660 95.055 62.705 ;
        RECT 97.705 62.660 98.355 62.705 ;
        RECT 94.465 62.520 98.720 62.660 ;
        RECT 94.465 62.475 94.755 62.520 ;
        RECT 97.705 62.475 98.355 62.520 ;
        RECT 92.970 62.120 93.290 62.380 ;
        RECT 98.580 62.320 98.720 62.520 ;
        RECT 100.330 62.460 100.650 62.720 ;
        RECT 103.180 62.380 103.320 62.815 ;
        RECT 111.920 62.705 112.060 62.860 ;
        RECT 111.845 62.475 112.135 62.705 ;
        RECT 112.380 62.660 112.520 63.540 ;
        RECT 113.635 63.540 118.935 63.680 ;
        RECT 113.635 63.495 113.925 63.540 ;
        RECT 115.525 63.495 115.815 63.540 ;
        RECT 118.645 63.495 118.935 63.540 ;
        RECT 119.740 63.540 122.640 63.680 ;
        RECT 142.280 63.540 143.430 63.680 ;
        RECT 112.750 62.800 113.070 63.060 ;
        RECT 113.230 63.000 113.520 63.045 ;
        RECT 115.065 63.000 115.355 63.045 ;
        RECT 118.645 63.000 118.935 63.045 ;
        RECT 119.740 63.020 119.880 63.540 ;
        RECT 121.030 63.340 121.350 63.400 ;
        RECT 142.280 63.340 142.420 63.540 ;
        RECT 143.110 63.480 143.430 63.540 ;
        RECT 146.420 63.340 146.560 63.820 ;
        RECT 121.030 63.200 142.420 63.340 ;
        RECT 121.030 63.140 121.350 63.200 ;
        RECT 142.280 63.045 142.420 63.200 ;
        RECT 143.200 63.200 146.560 63.340 ;
        RECT 143.200 63.045 143.340 63.200 ;
        RECT 113.230 62.860 118.935 63.000 ;
        RECT 113.230 62.815 113.520 62.860 ;
        RECT 115.065 62.815 115.355 62.860 ;
        RECT 118.645 62.815 118.935 62.860 ;
        RECT 113.670 62.660 113.990 62.720 ;
        RECT 112.380 62.520 113.990 62.660 ;
        RECT 102.645 62.320 102.935 62.365 ;
        RECT 98.580 62.180 102.935 62.320 ;
        RECT 102.645 62.135 102.935 62.180 ;
        RECT 103.090 62.120 103.410 62.380 ;
        RECT 105.850 62.120 106.170 62.380 ;
        RECT 107.230 62.120 107.550 62.380 ;
        RECT 107.690 62.320 108.010 62.380 ;
        RECT 109.545 62.320 109.835 62.365 ;
        RECT 107.690 62.180 109.835 62.320 ;
        RECT 111.920 62.320 112.060 62.475 ;
        RECT 113.670 62.460 113.990 62.520 ;
        RECT 114.130 62.460 114.450 62.720 ;
        RECT 119.725 62.705 120.015 63.020 ;
        RECT 124.725 62.815 125.015 63.045 ;
        RECT 126.565 63.000 126.855 63.045 ;
        RECT 126.180 62.860 126.855 63.000 ;
        RECT 116.425 62.660 117.075 62.705 ;
        RECT 119.725 62.660 120.315 62.705 ;
        RECT 124.800 62.660 124.940 62.815 ;
        RECT 116.425 62.520 120.315 62.660 ;
        RECT 116.425 62.475 117.075 62.520 ;
        RECT 120.025 62.475 120.315 62.520 ;
        RECT 121.580 62.520 124.940 62.660 ;
        RECT 121.580 62.365 121.720 62.520 ;
        RECT 126.180 62.380 126.320 62.860 ;
        RECT 126.565 62.815 126.855 62.860 ;
        RECT 142.205 62.815 142.495 63.045 ;
        RECT 143.125 62.815 143.415 63.045 ;
        RECT 146.330 63.000 146.650 63.060 ;
        RECT 147.265 63.000 147.555 63.045 ;
        RECT 146.330 62.860 147.555 63.000 ;
        RECT 146.330 62.800 146.650 62.860 ;
        RECT 147.265 62.815 147.555 62.860 ;
        RECT 121.505 62.320 121.795 62.365 ;
        RECT 111.920 62.180 121.795 62.320 ;
        RECT 107.690 62.120 108.010 62.180 ;
        RECT 109.545 62.135 109.835 62.180 ;
        RECT 121.505 62.135 121.795 62.180 ;
        RECT 121.950 62.120 122.270 62.380 ;
        RECT 126.090 62.120 126.410 62.380 ;
        RECT 142.650 62.120 142.970 62.380 ;
        RECT 88.980 61.500 152.240 61.980 ;
        RECT 55.390 56.715 56.290 57.505 ;
        RECT 88.980 56.540 89.460 61.500 ;
        RECT 92.970 61.300 93.290 61.360 ;
        RECT 95.730 61.300 96.050 61.360 ;
        RECT 100.330 61.300 100.650 61.360 ;
        RECT 101.725 61.300 102.015 61.345 ;
        RECT 92.970 61.160 99.410 61.300 ;
        RECT 92.970 61.100 93.290 61.160 ;
        RECT 95.730 61.100 96.050 61.160 ;
        RECT 97.585 60.960 97.875 61.005 ;
        RECT 99.270 60.960 99.410 61.160 ;
        RECT 100.330 61.160 102.015 61.300 ;
        RECT 100.330 61.100 100.650 61.160 ;
        RECT 101.725 61.115 102.015 61.160 ;
        RECT 102.185 61.300 102.475 61.345 ;
        RECT 103.550 61.300 103.870 61.360 ;
        RECT 102.185 61.160 103.870 61.300 ;
        RECT 102.185 61.115 102.475 61.160 ;
        RECT 103.550 61.100 103.870 61.160 ;
        RECT 107.230 61.100 107.550 61.360 ;
        RECT 114.130 61.100 114.450 61.360 ;
        RECT 115.985 61.300 116.275 61.345 ;
        RECT 121.950 61.300 122.270 61.360 ;
        RECT 115.985 61.160 122.270 61.300 ;
        RECT 115.985 61.115 116.275 61.160 ;
        RECT 121.950 61.100 122.270 61.160 ;
        RECT 138.050 61.100 138.370 61.360 ;
        RECT 146.330 61.100 146.650 61.360 ;
        RECT 103.105 60.960 103.395 61.005 ;
        RECT 105.405 60.960 105.695 61.005 ;
        RECT 97.585 60.820 98.720 60.960 ;
        RECT 99.270 60.820 100.560 60.960 ;
        RECT 97.585 60.775 97.875 60.820 ;
        RECT 97.125 60.435 97.415 60.665 ;
        RECT 97.200 59.940 97.340 60.435 ;
        RECT 98.030 60.420 98.350 60.680 ;
        RECT 98.580 60.665 98.720 60.820 ;
        RECT 98.505 60.435 98.795 60.665 ;
        RECT 99.410 60.420 99.730 60.680 ;
        RECT 99.870 60.420 100.190 60.680 ;
        RECT 100.420 60.665 100.560 60.820 ;
        RECT 103.105 60.820 105.695 60.960 ;
        RECT 107.320 60.960 107.460 61.100 ;
        RECT 115.510 60.960 115.830 61.020 ;
        RECT 117.365 60.960 117.655 61.005 ;
        RECT 107.320 60.820 107.920 60.960 ;
        RECT 103.105 60.775 103.395 60.820 ;
        RECT 105.405 60.775 105.695 60.820 ;
        RECT 100.345 60.620 100.635 60.665 ;
        RECT 102.170 60.620 102.490 60.680 ;
        RECT 100.345 60.480 102.490 60.620 ;
        RECT 100.345 60.435 100.635 60.480 ;
        RECT 102.170 60.420 102.490 60.480 ;
        RECT 104.930 60.620 105.250 60.680 ;
        RECT 106.325 60.620 106.615 60.665 ;
        RECT 106.770 60.620 107.090 60.680 ;
        RECT 104.930 60.480 107.090 60.620 ;
        RECT 104.930 60.420 105.250 60.480 ;
        RECT 106.325 60.435 106.615 60.480 ;
        RECT 106.770 60.420 107.090 60.480 ;
        RECT 107.230 60.420 107.550 60.680 ;
        RECT 107.780 60.665 107.920 60.820 ;
        RECT 115.510 60.820 117.655 60.960 ;
        RECT 115.510 60.760 115.830 60.820 ;
        RECT 117.365 60.775 117.655 60.820 ;
        RECT 107.705 60.435 107.995 60.665 ;
        RECT 113.670 60.620 113.990 60.680 ;
        RECT 115.065 60.620 115.355 60.665 ;
        RECT 113.670 60.480 115.355 60.620 ;
        RECT 100.790 60.280 101.110 60.340 ;
        RECT 107.780 60.280 107.920 60.435 ;
        RECT 113.670 60.420 113.990 60.480 ;
        RECT 115.065 60.435 115.355 60.480 ;
        RECT 116.445 60.620 116.735 60.665 ;
        RECT 127.010 60.620 127.330 60.680 ;
        RECT 116.445 60.480 127.330 60.620 ;
        RECT 116.445 60.435 116.735 60.480 ;
        RECT 99.270 60.140 107.920 60.280 ;
        RECT 115.140 60.280 115.280 60.435 ;
        RECT 127.010 60.420 127.330 60.480 ;
        RECT 138.140 60.280 138.280 61.100 ;
        RECT 146.420 60.960 146.560 61.100 ;
        RECT 147.265 60.960 147.555 61.005 ;
        RECT 146.420 60.820 147.555 60.960 ;
        RECT 147.265 60.775 147.555 60.820 ;
        RECT 145.870 60.420 146.190 60.680 ;
        RECT 115.140 60.140 138.280 60.280 ;
        RECT 99.270 59.940 99.410 60.140 ;
        RECT 100.790 60.080 101.110 60.140 ;
        RECT 150.010 60.080 150.330 60.340 ;
        RECT 97.200 59.800 99.410 59.940 ;
        RECT 104.945 59.940 105.235 59.985 ;
        RECT 105.850 59.940 106.170 60.000 ;
        RECT 104.945 59.800 106.170 59.940 ;
        RECT 104.945 59.755 105.235 59.800 ;
        RECT 105.850 59.740 106.170 59.800 ;
        RECT 146.345 59.940 146.635 59.985 ;
        RECT 146.345 59.800 147.940 59.940 ;
        RECT 146.345 59.755 146.635 59.800 ;
        RECT 147.800 59.660 147.940 59.800 ;
        RECT 96.650 59.600 96.970 59.660 ;
        RECT 99.410 59.600 99.730 59.660 ;
        RECT 103.105 59.600 103.395 59.645 ;
        RECT 108.610 59.600 108.930 59.660 ;
        RECT 96.650 59.460 108.930 59.600 ;
        RECT 96.650 59.400 96.970 59.460 ;
        RECT 99.410 59.400 99.730 59.460 ;
        RECT 103.105 59.415 103.395 59.460 ;
        RECT 108.610 59.400 108.930 59.460 ;
        RECT 123.790 59.400 124.110 59.660 ;
        RECT 147.710 59.400 148.030 59.660 ;
        RECT 152.900 59.260 153.380 64.220 ;
        RECT 91.060 58.780 153.380 59.260 ;
        RECT 96.650 58.380 96.970 58.640 ;
        RECT 98.505 58.580 98.795 58.625 ;
        RECT 99.870 58.580 100.190 58.640 ;
        RECT 98.505 58.440 100.190 58.580 ;
        RECT 98.505 58.395 98.795 58.440 ;
        RECT 96.740 57.945 96.880 58.380 ;
        RECT 96.665 57.715 96.955 57.945 ;
        RECT 97.570 57.360 97.890 57.620 ;
        RECT 98.045 57.560 98.335 57.605 ;
        RECT 98.580 57.560 98.720 58.395 ;
        RECT 99.870 58.380 100.190 58.440 ;
        RECT 100.790 58.380 101.110 58.640 ;
        RECT 107.230 58.380 107.550 58.640 ;
        RECT 110.910 58.580 111.230 58.640 ;
        RECT 113.225 58.580 113.515 58.625 ;
        RECT 110.910 58.440 113.515 58.580 ;
        RECT 110.910 58.380 111.230 58.440 ;
        RECT 113.225 58.395 113.515 58.440 ;
        RECT 150.010 58.380 150.330 58.640 ;
        RECT 107.320 57.900 107.460 58.380 ;
        RECT 142.155 58.240 142.445 58.285 ;
        RECT 144.045 58.240 144.335 58.285 ;
        RECT 147.165 58.240 147.455 58.285 ;
        RECT 142.155 58.100 147.455 58.240 ;
        RECT 142.155 58.055 142.445 58.100 ;
        RECT 144.045 58.055 144.335 58.100 ;
        RECT 147.165 58.055 147.455 58.100 ;
        RECT 99.500 57.760 107.460 57.900 ;
        RECT 131.150 57.900 131.470 57.960 ;
        RECT 132.085 57.900 132.375 57.945 ;
        RECT 131.150 57.760 132.375 57.900 ;
        RECT 98.045 57.420 98.720 57.560 ;
        RECT 98.950 57.560 99.270 57.620 ;
        RECT 99.500 57.605 99.640 57.760 ;
        RECT 131.150 57.700 131.470 57.760 ;
        RECT 132.085 57.715 132.375 57.760 ;
        RECT 142.650 57.700 142.970 57.960 ;
        RECT 99.425 57.560 99.715 57.605 ;
        RECT 100.330 57.560 100.650 57.620 ;
        RECT 101.725 57.560 102.015 57.605 ;
        RECT 98.950 57.420 99.925 57.560 ;
        RECT 100.330 57.420 102.015 57.560 ;
        RECT 98.045 57.375 98.335 57.420 ;
        RECT 98.950 57.360 99.270 57.420 ;
        RECT 99.425 57.375 99.715 57.420 ;
        RECT 100.330 57.360 100.650 57.420 ;
        RECT 101.725 57.375 102.015 57.420 ;
        RECT 102.170 57.360 102.490 57.620 ;
        RECT 120.570 57.560 120.890 57.620 ;
        RECT 123.790 57.560 124.110 57.620 ;
        RECT 120.570 57.420 124.110 57.560 ;
        RECT 120.570 57.360 120.890 57.420 ;
        RECT 123.790 57.360 124.110 57.420 ;
        RECT 126.090 57.360 126.410 57.620 ;
        RECT 126.565 57.560 126.855 57.605 ;
        RECT 127.930 57.560 128.250 57.620 ;
        RECT 126.565 57.420 128.250 57.560 ;
        RECT 126.565 57.375 126.855 57.420 ;
        RECT 127.930 57.360 128.250 57.420 ;
        RECT 133.925 57.560 134.215 57.605 ;
        RECT 135.290 57.560 135.610 57.620 ;
        RECT 133.925 57.420 135.610 57.560 ;
        RECT 133.925 57.375 134.215 57.420 ;
        RECT 135.290 57.360 135.610 57.420 ;
        RECT 141.270 57.360 141.590 57.620 ;
        RECT 141.750 57.560 142.040 57.605 ;
        RECT 143.585 57.560 143.875 57.605 ;
        RECT 147.165 57.560 147.455 57.605 ;
        RECT 141.750 57.420 147.455 57.560 ;
        RECT 141.750 57.375 142.040 57.420 ;
        RECT 143.585 57.375 143.875 57.420 ;
        RECT 147.165 57.375 147.455 57.420 ;
        RECT 97.110 57.220 97.430 57.280 ;
        RECT 99.040 57.220 99.180 57.360 ;
        RECT 126.180 57.220 126.320 57.360 ;
        RECT 97.110 57.080 99.180 57.220 ;
        RECT 118.360 57.080 126.320 57.220 ;
        RECT 97.110 57.020 97.430 57.080 ;
        RECT 118.360 56.940 118.500 57.080 ;
        RECT 130.230 57.020 130.550 57.280 ;
        RECT 131.165 57.220 131.455 57.265 ;
        RECT 136.210 57.220 136.530 57.280 ;
        RECT 131.165 57.080 136.530 57.220 ;
        RECT 131.165 57.035 131.455 57.080 ;
        RECT 136.210 57.020 136.530 57.080 ;
        RECT 144.945 57.220 145.595 57.265 ;
        RECT 147.710 57.220 148.030 57.280 ;
        RECT 148.245 57.265 148.535 57.580 ;
        RECT 148.245 57.220 148.835 57.265 ;
        RECT 144.945 57.080 148.835 57.220 ;
        RECT 144.945 57.035 145.595 57.080 ;
        RECT 147.710 57.020 148.030 57.080 ;
        RECT 148.545 57.035 148.835 57.080 ;
        RECT 96.650 56.680 96.970 56.940 ;
        RECT 118.270 56.680 118.590 56.940 ;
        RECT 125.630 56.680 125.950 56.940 ;
        RECT 127.470 56.680 127.790 56.940 ;
        RECT 133.005 56.880 133.295 56.925 ;
        RECT 133.450 56.880 133.770 56.940 ;
        RECT 133.005 56.740 133.770 56.880 ;
        RECT 133.005 56.695 133.295 56.740 ;
        RECT 133.450 56.680 133.770 56.740 ;
        RECT 88.980 56.060 152.240 56.540 ;
        RECT 6.020 50.910 6.380 51.050 ;
        RECT 25.005 50.885 27.255 51.165 ;
        RECT 6.080 44.445 6.330 46.550 ;
        RECT 6.080 41.290 6.330 43.395 ;
        RECT 26.975 37.600 27.255 50.885 ;
        RECT 5.965 37.320 27.255 37.600 ;
        RECT 88.980 51.100 89.460 56.060 ;
        RECT 97.570 55.860 97.890 55.920 ;
        RECT 98.965 55.860 99.255 55.905 ;
        RECT 97.570 55.720 99.255 55.860 ;
        RECT 97.570 55.660 97.890 55.720 ;
        RECT 98.965 55.675 99.255 55.720 ;
        RECT 115.065 55.860 115.355 55.905 ;
        RECT 115.065 55.720 116.660 55.860 ;
        RECT 115.065 55.675 115.355 55.720 ;
        RECT 114.145 55.520 114.435 55.565 ;
        RECT 114.145 55.380 115.280 55.520 ;
        RECT 114.145 55.335 114.435 55.380 ;
        RECT 115.140 55.240 115.280 55.380 ;
        RECT 98.505 55.180 98.795 55.225 ;
        RECT 98.950 55.180 99.270 55.240 ;
        RECT 98.505 55.040 99.270 55.180 ;
        RECT 98.505 54.995 98.795 55.040 ;
        RECT 98.950 54.980 99.270 55.040 ;
        RECT 99.425 55.180 99.715 55.225 ;
        RECT 100.330 55.180 100.650 55.240 ;
        RECT 99.425 55.040 100.650 55.180 ;
        RECT 99.425 54.995 99.715 55.040 ;
        RECT 100.330 54.980 100.650 55.040 ;
        RECT 103.090 54.980 103.410 55.240 ;
        RECT 115.050 54.980 115.370 55.240 ;
        RECT 116.520 55.225 116.660 55.720 ;
        RECT 127.470 55.660 127.790 55.920 ;
        RECT 131.700 55.720 141.500 55.860 ;
        RECT 123.445 55.520 123.735 55.565 ;
        RECT 125.630 55.520 125.950 55.580 ;
        RECT 126.685 55.520 127.335 55.565 ;
        RECT 123.445 55.380 127.335 55.520 ;
        RECT 127.560 55.520 127.700 55.660 ;
        RECT 129.325 55.520 129.615 55.565 ;
        RECT 127.560 55.380 129.615 55.520 ;
        RECT 123.445 55.335 124.035 55.380 ;
        RECT 116.445 54.995 116.735 55.225 ;
        RECT 118.270 54.980 118.590 55.240 ;
        RECT 123.745 55.020 124.035 55.335 ;
        RECT 125.630 55.320 125.950 55.380 ;
        RECT 126.685 55.335 127.335 55.380 ;
        RECT 129.325 55.335 129.615 55.380 ;
        RECT 124.825 55.180 125.115 55.225 ;
        RECT 128.405 55.180 128.695 55.225 ;
        RECT 130.240 55.180 130.530 55.225 ;
        RECT 124.825 55.040 130.530 55.180 ;
        RECT 124.825 54.995 125.115 55.040 ;
        RECT 128.405 54.995 128.695 55.040 ;
        RECT 130.240 54.995 130.530 55.040 ;
        RECT 130.690 55.180 131.010 55.240 ;
        RECT 131.700 55.225 131.840 55.720 ;
        RECT 141.360 55.580 141.500 55.720 ;
        RECT 133.005 55.520 133.295 55.565 ;
        RECT 133.450 55.520 133.770 55.580 ;
        RECT 133.005 55.380 133.770 55.520 ;
        RECT 133.005 55.335 133.295 55.380 ;
        RECT 133.450 55.320 133.770 55.380 ;
        RECT 135.285 55.520 135.935 55.565 ;
        RECT 138.885 55.520 139.175 55.565 ;
        RECT 135.285 55.380 139.175 55.520 ;
        RECT 135.285 55.335 135.935 55.380 ;
        RECT 138.585 55.335 139.175 55.380 ;
        RECT 131.625 55.180 131.915 55.225 ;
        RECT 130.690 55.040 131.915 55.180 ;
        RECT 130.690 54.980 131.010 55.040 ;
        RECT 131.625 54.995 131.915 55.040 ;
        RECT 132.090 55.180 132.380 55.225 ;
        RECT 133.925 55.180 134.215 55.225 ;
        RECT 137.505 55.180 137.795 55.225 ;
        RECT 132.090 55.040 137.795 55.180 ;
        RECT 132.090 54.995 132.380 55.040 ;
        RECT 133.925 54.995 134.215 55.040 ;
        RECT 137.505 54.995 137.795 55.040 ;
        RECT 138.585 55.020 138.875 55.335 ;
        RECT 141.270 55.320 141.590 55.580 ;
        RECT 141.745 55.180 142.035 55.225 ;
        RECT 145.870 55.180 146.190 55.240 ;
        RECT 146.345 55.180 146.635 55.225 ;
        RECT 141.745 55.040 146.635 55.180 ;
        RECT 103.180 54.840 103.320 54.980 ;
        RECT 118.360 54.840 118.500 54.980 ;
        RECT 103.180 54.700 118.500 54.840 ;
        RECT 138.600 54.840 138.740 55.020 ;
        RECT 141.745 54.995 142.035 55.040 ;
        RECT 141.285 54.840 141.575 54.885 ;
        RECT 138.600 54.700 141.575 54.840 ;
        RECT 141.820 54.840 141.960 54.995 ;
        RECT 145.870 54.980 146.190 55.040 ;
        RECT 146.345 54.995 146.635 55.040 ;
        RECT 142.650 54.840 142.970 54.900 ;
        RECT 141.820 54.700 142.970 54.840 ;
        RECT 141.285 54.655 141.575 54.700 ;
        RECT 142.650 54.640 142.970 54.700 ;
        RECT 110.450 54.500 110.770 54.560 ;
        RECT 112.305 54.500 112.595 54.545 ;
        RECT 124.825 54.500 125.115 54.545 ;
        RECT 127.945 54.500 128.235 54.545 ;
        RECT 129.835 54.500 130.125 54.545 ;
        RECT 110.450 54.360 112.595 54.500 ;
        RECT 110.450 54.300 110.770 54.360 ;
        RECT 112.305 54.315 112.595 54.360 ;
        RECT 115.140 54.360 118.500 54.500 ;
        RECT 108.610 54.160 108.930 54.220 ;
        RECT 114.145 54.160 114.435 54.205 ;
        RECT 115.140 54.160 115.280 54.360 ;
        RECT 118.360 54.220 118.500 54.360 ;
        RECT 124.825 54.360 130.125 54.500 ;
        RECT 124.825 54.315 125.115 54.360 ;
        RECT 127.945 54.315 128.235 54.360 ;
        RECT 129.835 54.315 130.125 54.360 ;
        RECT 132.495 54.500 132.785 54.545 ;
        RECT 134.385 54.500 134.675 54.545 ;
        RECT 137.505 54.500 137.795 54.545 ;
        RECT 132.495 54.360 137.795 54.500 ;
        RECT 132.495 54.315 132.785 54.360 ;
        RECT 134.385 54.315 134.675 54.360 ;
        RECT 137.505 54.315 137.795 54.360 ;
        RECT 108.610 54.020 115.280 54.160 ;
        RECT 108.610 53.960 108.930 54.020 ;
        RECT 114.145 53.975 114.435 54.020 ;
        RECT 115.510 53.960 115.830 54.220 ;
        RECT 118.270 53.960 118.590 54.220 ;
        RECT 118.745 54.160 119.035 54.205 ;
        RECT 120.110 54.160 120.430 54.220 ;
        RECT 118.745 54.020 120.430 54.160 ;
        RECT 118.745 53.975 119.035 54.020 ;
        RECT 120.110 53.960 120.430 54.020 ;
        RECT 121.950 53.960 122.270 54.220 ;
        RECT 136.210 54.160 136.530 54.220 ;
        RECT 140.365 54.160 140.655 54.205 ;
        RECT 136.210 54.020 140.655 54.160 ;
        RECT 136.210 53.960 136.530 54.020 ;
        RECT 140.365 53.975 140.655 54.020 ;
        RECT 146.805 54.160 147.095 54.205 ;
        RECT 147.710 54.160 148.030 54.220 ;
        RECT 146.805 54.020 148.030 54.160 ;
        RECT 146.805 53.975 147.095 54.020 ;
        RECT 147.710 53.960 148.030 54.020 ;
        RECT 152.900 53.820 153.380 58.780 ;
        RECT 91.060 53.340 153.380 53.820 ;
        RECT 93.840 53.140 94.130 53.185 ;
        RECT 96.650 53.140 96.970 53.200 ;
        RECT 93.840 53.000 96.970 53.140 ;
        RECT 93.840 52.955 94.130 53.000 ;
        RECT 96.650 52.940 96.970 53.000 ;
        RECT 114.540 53.140 114.830 53.185 ;
        RECT 115.510 53.140 115.830 53.200 ;
        RECT 114.540 53.000 115.830 53.140 ;
        RECT 114.540 52.955 114.830 53.000 ;
        RECT 115.510 52.940 115.830 53.000 ;
        RECT 118.270 53.140 118.590 53.200 ;
        RECT 127.485 53.140 127.775 53.185 ;
        RECT 118.270 53.000 127.775 53.140 ;
        RECT 118.270 52.940 118.590 53.000 ;
        RECT 127.485 52.955 127.775 53.000 ;
        RECT 127.930 53.140 128.250 53.200 ;
        RECT 128.405 53.140 128.695 53.185 ;
        RECT 132.085 53.140 132.375 53.185 ;
        RECT 127.930 53.000 128.695 53.140 ;
        RECT 93.395 52.800 93.685 52.845 ;
        RECT 95.285 52.800 95.575 52.845 ;
        RECT 98.405 52.800 98.695 52.845 ;
        RECT 93.395 52.660 98.695 52.800 ;
        RECT 93.395 52.615 93.685 52.660 ;
        RECT 95.285 52.615 95.575 52.660 ;
        RECT 98.405 52.615 98.695 52.660 ;
        RECT 114.095 52.800 114.385 52.845 ;
        RECT 115.985 52.800 116.275 52.845 ;
        RECT 119.105 52.800 119.395 52.845 ;
        RECT 114.095 52.660 119.395 52.800 ;
        RECT 127.560 52.800 127.700 52.955 ;
        RECT 127.930 52.940 128.250 53.000 ;
        RECT 128.405 52.955 128.695 53.000 ;
        RECT 128.940 53.000 132.375 53.140 ;
        RECT 128.940 52.800 129.080 53.000 ;
        RECT 132.085 52.955 132.375 53.000 ;
        RECT 133.450 53.140 133.770 53.200 ;
        RECT 135.305 53.140 135.595 53.185 ;
        RECT 133.450 53.000 135.595 53.140 ;
        RECT 127.560 52.660 129.080 52.800 ;
        RECT 114.095 52.615 114.385 52.660 ;
        RECT 115.985 52.615 116.275 52.660 ;
        RECT 119.105 52.615 119.395 52.660 ;
        RECT 131.165 52.615 131.455 52.845 ;
        RECT 132.160 52.800 132.300 52.955 ;
        RECT 133.450 52.940 133.770 53.000 ;
        RECT 135.305 52.955 135.595 53.000 ;
        RECT 138.525 53.140 138.815 53.185 ;
        RECT 140.350 53.140 140.670 53.200 ;
        RECT 138.525 53.000 140.670 53.140 ;
        RECT 138.525 52.955 138.815 53.000 ;
        RECT 138.600 52.800 138.740 52.955 ;
        RECT 140.350 52.940 140.670 53.000 ;
        RECT 132.160 52.660 138.740 52.800 ;
        RECT 142.155 52.800 142.445 52.845 ;
        RECT 144.045 52.800 144.335 52.845 ;
        RECT 147.165 52.800 147.455 52.845 ;
        RECT 142.155 52.660 147.455 52.800 ;
        RECT 142.155 52.615 142.445 52.660 ;
        RECT 144.045 52.615 144.335 52.660 ;
        RECT 147.165 52.615 147.455 52.660 ;
        RECT 106.310 52.460 106.630 52.520 ;
        RECT 110.910 52.460 111.230 52.520 ;
        RECT 112.750 52.460 113.070 52.520 ;
        RECT 113.225 52.460 113.515 52.505 ;
        RECT 131.240 52.460 131.380 52.615 ;
        RECT 135.290 52.460 135.610 52.520 ;
        RECT 106.310 52.320 110.680 52.460 ;
        RECT 106.310 52.260 106.630 52.320 ;
        RECT 92.510 51.920 92.830 52.180 ;
        RECT 92.990 52.120 93.280 52.165 ;
        RECT 94.825 52.120 95.115 52.165 ;
        RECT 98.405 52.120 98.695 52.165 ;
        RECT 92.990 51.980 98.695 52.120 ;
        RECT 92.990 51.935 93.280 51.980 ;
        RECT 94.825 51.935 95.115 51.980 ;
        RECT 98.405 51.935 98.695 51.980 ;
        RECT 99.485 51.825 99.775 52.140 ;
        RECT 100.790 52.120 101.110 52.180 ;
        RECT 102.645 52.120 102.935 52.165 ;
        RECT 103.090 52.120 103.410 52.180 ;
        RECT 100.790 51.980 103.410 52.120 ;
        RECT 100.790 51.920 101.110 51.980 ;
        RECT 102.645 51.935 102.935 51.980 ;
        RECT 103.090 51.920 103.410 51.980 ;
        RECT 109.990 51.920 110.310 52.180 ;
        RECT 110.540 52.120 110.680 52.320 ;
        RECT 110.910 52.320 130.920 52.460 ;
        RECT 131.240 52.320 135.610 52.460 ;
        RECT 110.910 52.260 111.230 52.320 ;
        RECT 112.750 52.260 113.070 52.320 ;
        RECT 113.225 52.275 113.515 52.320 ;
        RECT 130.780 52.180 130.920 52.320 ;
        RECT 135.290 52.260 135.610 52.320 ;
        RECT 137.590 52.460 137.910 52.520 ;
        RECT 150.025 52.460 150.315 52.505 ;
        RECT 137.590 52.320 150.315 52.460 ;
        RECT 137.590 52.260 137.910 52.320 ;
        RECT 150.025 52.275 150.315 52.320 ;
        RECT 111.370 52.120 111.690 52.180 ;
        RECT 110.540 51.980 111.690 52.120 ;
        RECT 111.370 51.920 111.690 51.980 ;
        RECT 113.690 52.120 113.980 52.165 ;
        RECT 115.525 52.120 115.815 52.165 ;
        RECT 119.105 52.120 119.395 52.165 ;
        RECT 113.690 51.980 119.395 52.120 ;
        RECT 113.690 51.935 113.980 51.980 ;
        RECT 115.525 51.935 115.815 51.980 ;
        RECT 119.105 51.935 119.395 51.980 ;
        RECT 120.110 52.140 120.430 52.180 ;
        RECT 120.110 51.920 120.475 52.140 ;
        RECT 121.950 52.120 122.270 52.180 ;
        RECT 123.345 52.120 123.635 52.165 ;
        RECT 121.950 51.980 123.635 52.120 ;
        RECT 121.950 51.920 122.270 51.980 ;
        RECT 123.345 51.935 123.635 51.980 ;
        RECT 124.265 51.935 124.555 52.165 ;
        RECT 125.185 52.120 125.475 52.165 ;
        RECT 125.645 52.120 125.935 52.165 ;
        RECT 130.230 52.120 130.550 52.180 ;
        RECT 125.185 51.980 130.550 52.120 ;
        RECT 125.185 51.935 125.475 51.980 ;
        RECT 125.645 51.935 125.935 51.980 ;
        RECT 96.185 51.780 96.835 51.825 ;
        RECT 99.485 51.780 100.075 51.825 ;
        RECT 102.185 51.780 102.475 51.825 ;
        RECT 96.185 51.640 102.475 51.780 ;
        RECT 96.185 51.595 96.835 51.640 ;
        RECT 99.785 51.595 100.075 51.640 ;
        RECT 102.185 51.595 102.475 51.640 ;
        RECT 104.010 51.780 104.330 51.840 ;
        RECT 106.325 51.780 106.615 51.825 ;
        RECT 104.010 51.640 106.615 51.780 ;
        RECT 104.010 51.580 104.330 51.640 ;
        RECT 106.325 51.595 106.615 51.640 ;
        RECT 106.770 51.780 107.090 51.840 ;
        RECT 107.245 51.780 107.535 51.825 ;
        RECT 106.770 51.640 107.535 51.780 ;
        RECT 106.770 51.580 107.090 51.640 ;
        RECT 107.245 51.595 107.535 51.640 ;
        RECT 107.690 51.780 108.010 51.840 ;
        RECT 110.925 51.780 111.215 51.825 ;
        RECT 107.690 51.640 111.215 51.780 ;
        RECT 107.690 51.580 108.010 51.640 ;
        RECT 110.925 51.595 111.215 51.640 ;
        RECT 111.845 51.780 112.135 51.825 ;
        RECT 112.290 51.780 112.610 51.840 ;
        RECT 111.845 51.640 112.610 51.780 ;
        RECT 111.845 51.595 112.135 51.640 ;
        RECT 112.290 51.580 112.610 51.640 ;
        RECT 112.765 51.780 113.055 51.825 ;
        RECT 115.050 51.780 115.370 51.840 ;
        RECT 120.185 51.825 120.475 51.920 ;
        RECT 112.765 51.640 115.370 51.780 ;
        RECT 112.765 51.595 113.055 51.640 ;
        RECT 115.050 51.580 115.370 51.640 ;
        RECT 116.885 51.780 117.535 51.825 ;
        RECT 120.185 51.780 120.775 51.825 ;
        RECT 116.885 51.640 120.775 51.780 ;
        RECT 116.885 51.595 117.535 51.640 ;
        RECT 120.485 51.595 120.775 51.640 ;
        RECT 121.490 51.780 121.810 51.840 ;
        RECT 124.340 51.780 124.480 51.935 ;
        RECT 130.230 51.920 130.550 51.980 ;
        RECT 130.690 51.920 131.010 52.180 ;
        RECT 131.150 52.120 131.470 52.180 ;
        RECT 131.150 51.980 132.300 52.120 ;
        RECT 131.150 51.920 131.470 51.980 ;
        RECT 132.160 51.825 132.300 51.980 ;
        RECT 133.925 51.935 134.215 52.165 ;
        RECT 121.490 51.640 124.480 51.780 ;
        RECT 121.490 51.580 121.810 51.640 ;
        RECT 132.085 51.595 132.375 51.825 ;
        RECT 100.330 51.440 100.650 51.500 ;
        RECT 101.265 51.440 101.555 51.485 ;
        RECT 100.330 51.300 101.555 51.440 ;
        RECT 100.330 51.240 100.650 51.300 ;
        RECT 101.265 51.255 101.555 51.300 ;
        RECT 108.150 51.240 108.470 51.500 ;
        RECT 109.070 51.240 109.390 51.500 ;
        RECT 112.380 51.440 112.520 51.580 ;
        RECT 121.965 51.440 122.255 51.485 ;
        RECT 122.410 51.440 122.730 51.500 ;
        RECT 112.380 51.300 122.730 51.440 ;
        RECT 121.965 51.255 122.255 51.300 ;
        RECT 122.410 51.240 122.730 51.300 ;
        RECT 127.470 51.240 127.790 51.500 ;
        RECT 134.000 51.440 134.140 51.935 ;
        RECT 134.370 51.920 134.690 52.180 ;
        RECT 134.830 52.120 135.150 52.180 ;
        RECT 136.685 52.120 136.975 52.165 ;
        RECT 139.905 52.120 140.195 52.165 ;
        RECT 134.830 51.980 136.975 52.120 ;
        RECT 134.830 51.920 135.150 51.980 ;
        RECT 136.685 51.935 136.975 51.980 ;
        RECT 139.520 51.980 140.195 52.120 ;
        RECT 134.460 51.780 134.600 51.920 ;
        RECT 134.460 51.640 135.060 51.780 ;
        RECT 134.370 51.440 134.690 51.500 ;
        RECT 134.000 51.300 134.690 51.440 ;
        RECT 134.920 51.440 135.060 51.640 ;
        RECT 136.210 51.580 136.530 51.840 ;
        RECT 135.225 51.440 135.515 51.485 ;
        RECT 134.920 51.300 135.515 51.440 ;
        RECT 134.370 51.240 134.690 51.300 ;
        RECT 135.225 51.255 135.515 51.300 ;
        RECT 138.510 51.240 138.830 51.500 ;
        RECT 139.520 51.485 139.660 51.980 ;
        RECT 139.905 51.935 140.195 51.980 ;
        RECT 141.270 51.920 141.590 52.180 ;
        RECT 141.750 52.120 142.040 52.165 ;
        RECT 143.585 52.120 143.875 52.165 ;
        RECT 147.165 52.120 147.455 52.165 ;
        RECT 141.750 51.980 147.455 52.120 ;
        RECT 141.750 51.935 142.040 51.980 ;
        RECT 143.585 51.935 143.875 51.980 ;
        RECT 147.165 51.935 147.455 51.980 ;
        RECT 142.665 51.780 142.955 51.825 ;
        RECT 140.900 51.640 142.955 51.780 ;
        RECT 140.900 51.485 141.040 51.640 ;
        RECT 142.665 51.595 142.955 51.640 ;
        RECT 144.945 51.780 145.595 51.825 ;
        RECT 147.710 51.780 148.030 51.840 ;
        RECT 148.245 51.825 148.535 52.140 ;
        RECT 148.245 51.780 148.835 51.825 ;
        RECT 144.945 51.640 148.835 51.780 ;
        RECT 144.945 51.595 145.595 51.640 ;
        RECT 147.710 51.580 148.030 51.640 ;
        RECT 148.545 51.595 148.835 51.640 ;
        RECT 139.445 51.255 139.735 51.485 ;
        RECT 140.825 51.255 141.115 51.485 ;
        RECT 88.980 50.620 152.240 51.100 ;
        RECT 88.980 45.660 89.460 50.620 ;
        RECT 104.945 50.420 105.235 50.465 ;
        RECT 107.690 50.420 108.010 50.480 ;
        RECT 104.945 50.280 108.010 50.420 ;
        RECT 104.945 50.235 105.235 50.280 ;
        RECT 107.690 50.220 108.010 50.280 ;
        RECT 109.070 50.220 109.390 50.480 ;
        RECT 110.450 50.420 110.770 50.480 ;
        RECT 121.490 50.420 121.810 50.480 ;
        RECT 110.450 50.280 121.810 50.420 ;
        RECT 110.450 50.220 110.770 50.280 ;
        RECT 121.490 50.220 121.810 50.280 ;
        RECT 127.470 50.420 127.790 50.480 ;
        RECT 128.405 50.420 128.695 50.465 ;
        RECT 127.470 50.280 128.695 50.420 ;
        RECT 127.470 50.220 127.790 50.280 ;
        RECT 128.405 50.235 128.695 50.280 ;
        RECT 128.850 50.420 129.170 50.480 ;
        RECT 133.910 50.420 134.230 50.480 ;
        RECT 128.850 50.280 134.230 50.420 ;
        RECT 128.850 50.220 129.170 50.280 ;
        RECT 133.910 50.220 134.230 50.280 ;
        RECT 134.370 50.420 134.690 50.480 ;
        RECT 134.370 50.280 135.520 50.420 ;
        RECT 134.370 50.220 134.690 50.280 ;
        RECT 92.510 50.080 92.830 50.140 ;
        RECT 92.510 49.940 102.860 50.080 ;
        RECT 92.510 49.880 92.830 49.940 ;
        RECT 98.505 49.740 98.795 49.785 ;
        RECT 99.885 49.740 100.175 49.785 ;
        RECT 101.250 49.740 101.570 49.800 ;
        RECT 98.505 49.600 99.410 49.740 ;
        RECT 98.505 49.555 98.795 49.600 ;
        RECT 97.110 49.200 97.430 49.460 ;
        RECT 99.270 49.400 99.410 49.600 ;
        RECT 99.885 49.600 101.570 49.740 ;
        RECT 99.885 49.555 100.175 49.600 ;
        RECT 101.250 49.540 101.570 49.600 ;
        RECT 100.790 49.400 101.110 49.460 ;
        RECT 99.270 49.260 101.110 49.400 ;
        RECT 100.790 49.200 101.110 49.260 ;
        RECT 97.200 49.060 97.340 49.200 ;
        RECT 101.340 49.060 101.480 49.540 ;
        RECT 102.185 49.215 102.475 49.445 ;
        RECT 102.720 49.400 102.860 49.940 ;
        RECT 105.635 49.910 105.925 49.955 ;
        RECT 103.105 49.740 103.395 49.785 ;
        RECT 105.635 49.740 106.000 49.910 ;
        RECT 106.770 49.880 107.090 50.140 ;
        RECT 108.625 50.080 108.915 50.125 ;
        RECT 109.160 50.080 109.300 50.220 ;
        RECT 108.625 49.940 109.300 50.080 ;
        RECT 110.905 50.080 111.555 50.125 ;
        RECT 114.505 50.080 114.795 50.125 ;
        RECT 115.050 50.080 115.370 50.140 ;
        RECT 110.905 49.940 115.370 50.080 ;
        RECT 108.625 49.895 108.915 49.940 ;
        RECT 110.905 49.895 111.555 49.940 ;
        RECT 114.205 49.895 114.795 49.940 ;
        RECT 107.245 49.740 107.535 49.785 ;
        RECT 103.105 49.600 106.000 49.740 ;
        RECT 103.105 49.555 103.395 49.600 ;
        RECT 105.860 49.460 106.000 49.600 ;
        RECT 106.400 49.600 107.535 49.740 ;
        RECT 102.720 49.260 103.320 49.400 ;
        RECT 97.200 48.920 101.480 49.060 ;
        RECT 102.260 49.060 102.400 49.215 ;
        RECT 103.180 49.060 103.320 49.260 ;
        RECT 104.010 49.200 104.330 49.460 ;
        RECT 105.850 49.200 106.170 49.460 ;
        RECT 106.400 49.060 106.540 49.600 ;
        RECT 107.245 49.555 107.535 49.600 ;
        RECT 107.710 49.740 108.000 49.785 ;
        RECT 109.545 49.740 109.835 49.785 ;
        RECT 113.125 49.740 113.415 49.785 ;
        RECT 107.710 49.600 113.415 49.740 ;
        RECT 107.710 49.555 108.000 49.600 ;
        RECT 109.545 49.555 109.835 49.600 ;
        RECT 113.125 49.555 113.415 49.600 ;
        RECT 114.205 49.580 114.495 49.895 ;
        RECT 115.050 49.880 115.370 49.940 ;
        RECT 121.580 49.740 121.720 50.220 ;
        RECT 121.950 50.080 122.270 50.140 ;
        RECT 131.150 50.080 131.470 50.140 ;
        RECT 133.005 50.080 133.295 50.125 ;
        RECT 121.950 49.940 128.620 50.080 ;
        RECT 121.950 49.880 122.270 49.940 ;
        RECT 127.560 49.785 127.700 49.940 ;
        RECT 126.565 49.740 126.855 49.785 ;
        RECT 121.580 49.600 126.855 49.740 ;
        RECT 126.565 49.555 126.855 49.600 ;
        RECT 127.485 49.555 127.775 49.785 ;
        RECT 128.480 49.740 128.620 49.940 ;
        RECT 131.150 49.940 134.600 50.080 ;
        RECT 131.150 49.880 131.470 49.940 ;
        RECT 133.005 49.895 133.295 49.940 ;
        RECT 133.450 49.740 133.770 49.800 ;
        RECT 128.480 49.600 133.770 49.740 ;
        RECT 134.460 49.740 134.600 49.940 ;
        RECT 134.830 49.880 135.150 50.140 ;
        RECT 135.380 50.125 135.520 50.280 ;
        RECT 135.750 50.220 136.070 50.480 ;
        RECT 137.145 50.420 137.435 50.465 ;
        RECT 138.510 50.420 138.830 50.480 ;
        RECT 137.145 50.280 138.830 50.420 ;
        RECT 137.145 50.235 137.435 50.280 ;
        RECT 138.510 50.220 138.830 50.280 ;
        RECT 135.305 49.895 135.595 50.125 ;
        RECT 135.840 49.740 135.980 50.220 ;
        RECT 136.225 50.080 136.515 50.125 ;
        RECT 137.590 50.080 137.910 50.140 ;
        RECT 136.225 49.940 137.910 50.080 ;
        RECT 136.225 49.895 136.515 49.940 ;
        RECT 134.460 49.600 135.980 49.740 ;
        RECT 106.770 49.400 107.090 49.460 ;
        RECT 111.830 49.400 112.150 49.460 ;
        RECT 115.985 49.400 116.275 49.445 ;
        RECT 106.770 49.260 116.275 49.400 ;
        RECT 126.640 49.400 126.780 49.555 ;
        RECT 133.450 49.540 133.770 49.600 ;
        RECT 128.850 49.400 129.170 49.460 ;
        RECT 126.640 49.260 129.170 49.400 ;
        RECT 106.770 49.200 107.090 49.260 ;
        RECT 111.830 49.200 112.150 49.260 ;
        RECT 115.985 49.215 116.275 49.260 ;
        RECT 128.850 49.200 129.170 49.260 ;
        RECT 132.085 49.400 132.375 49.445 ;
        RECT 134.370 49.400 134.690 49.460 ;
        RECT 136.300 49.400 136.440 49.895 ;
        RECT 137.590 49.880 137.910 49.940 ;
        RECT 145.410 49.740 145.730 49.800 ;
        RECT 149.105 49.740 149.395 49.785 ;
        RECT 145.410 49.600 149.395 49.740 ;
        RECT 145.410 49.540 145.730 49.600 ;
        RECT 149.105 49.555 149.395 49.600 ;
        RECT 132.085 49.260 136.440 49.400 ;
        RECT 132.085 49.215 132.375 49.260 ;
        RECT 134.370 49.200 134.690 49.260 ;
        RECT 150.470 49.200 150.790 49.460 ;
        RECT 102.260 48.920 102.860 49.060 ;
        RECT 103.180 48.920 106.540 49.060 ;
        RECT 96.190 48.720 96.510 48.780 ;
        RECT 97.585 48.720 97.875 48.765 ;
        RECT 96.190 48.580 97.875 48.720 ;
        RECT 96.190 48.520 96.510 48.580 ;
        RECT 97.585 48.535 97.875 48.580 ;
        RECT 99.425 48.720 99.715 48.765 ;
        RECT 99.870 48.720 100.190 48.780 ;
        RECT 99.425 48.580 100.190 48.720 ;
        RECT 102.720 48.720 102.860 48.920 ;
        RECT 105.390 48.720 105.710 48.780 ;
        RECT 105.865 48.720 106.155 48.765 ;
        RECT 102.720 48.580 106.155 48.720 ;
        RECT 106.400 48.720 106.540 48.920 ;
        RECT 108.115 49.060 108.405 49.105 ;
        RECT 110.005 49.060 110.295 49.105 ;
        RECT 113.125 49.060 113.415 49.105 ;
        RECT 108.115 48.920 113.415 49.060 ;
        RECT 108.115 48.875 108.405 48.920 ;
        RECT 110.005 48.875 110.295 48.920 ;
        RECT 113.125 48.875 113.415 48.920 ;
        RECT 110.910 48.720 111.230 48.780 ;
        RECT 106.400 48.580 111.230 48.720 ;
        RECT 99.425 48.535 99.715 48.580 ;
        RECT 99.870 48.520 100.190 48.580 ;
        RECT 105.390 48.520 105.710 48.580 ;
        RECT 105.865 48.535 106.155 48.580 ;
        RECT 110.910 48.520 111.230 48.580 ;
        RECT 152.900 48.380 153.380 53.340 ;
        RECT 91.060 47.900 153.380 48.380 ;
        RECT 92.510 47.500 92.830 47.760 ;
        RECT 107.230 47.500 107.550 47.760 ;
        RECT 107.690 47.500 108.010 47.760 ;
        RECT 108.150 47.500 108.470 47.760 ;
        RECT 109.990 47.500 110.310 47.760 ;
        RECT 110.910 47.500 111.230 47.760 ;
        RECT 111.370 47.700 111.690 47.760 ;
        RECT 117.825 47.700 118.115 47.745 ;
        RECT 120.110 47.700 120.430 47.760 ;
        RECT 111.370 47.560 120.430 47.700 ;
        RECT 111.370 47.500 111.690 47.560 ;
        RECT 117.825 47.515 118.115 47.560 ;
        RECT 120.110 47.500 120.430 47.560 ;
        RECT 92.600 47.020 92.740 47.500 ;
        RECT 93.855 47.360 94.145 47.405 ;
        RECT 95.745 47.360 96.035 47.405 ;
        RECT 98.865 47.360 99.155 47.405 ;
        RECT 93.855 47.220 99.155 47.360 ;
        RECT 93.855 47.175 94.145 47.220 ;
        RECT 95.745 47.175 96.035 47.220 ;
        RECT 98.865 47.175 99.155 47.220 ;
        RECT 105.405 47.360 105.695 47.405 ;
        RECT 107.780 47.360 107.920 47.500 ;
        RECT 105.405 47.220 107.920 47.360 ;
        RECT 105.405 47.175 105.695 47.220 ;
        RECT 92.985 47.020 93.275 47.065 ;
        RECT 92.600 46.880 93.275 47.020 ;
        RECT 92.985 46.835 93.275 46.880 ;
        RECT 94.365 47.020 94.655 47.065 ;
        RECT 96.190 47.020 96.510 47.080 ;
        RECT 94.365 46.880 96.510 47.020 ;
        RECT 94.365 46.835 94.655 46.880 ;
        RECT 96.190 46.820 96.510 46.880 ;
        RECT 93.450 46.680 93.740 46.725 ;
        RECT 95.285 46.680 95.575 46.725 ;
        RECT 98.865 46.680 99.155 46.725 ;
        RECT 93.450 46.540 99.155 46.680 ;
        RECT 93.450 46.495 93.740 46.540 ;
        RECT 95.285 46.495 95.575 46.540 ;
        RECT 98.865 46.495 99.155 46.540 ;
        RECT 99.870 46.700 100.190 46.740 ;
        RECT 99.870 46.480 100.235 46.700 ;
        RECT 99.945 46.385 100.235 46.480 ;
        RECT 96.645 46.340 97.295 46.385 ;
        RECT 99.945 46.340 100.535 46.385 ;
        RECT 96.645 46.200 100.535 46.340 ;
        RECT 96.645 46.155 97.295 46.200 ;
        RECT 100.245 46.155 100.535 46.200 ;
        RECT 107.245 46.340 107.535 46.385 ;
        RECT 108.240 46.340 108.380 47.500 ;
        RECT 107.245 46.200 108.380 46.340 ;
        RECT 107.245 46.155 107.535 46.200 ;
        RECT 101.725 46.000 102.015 46.045 ;
        RECT 105.390 46.000 105.710 46.060 ;
        RECT 101.725 45.860 105.710 46.000 ;
        RECT 101.725 45.815 102.015 45.860 ;
        RECT 105.390 45.800 105.710 45.860 ;
        RECT 108.165 46.000 108.455 46.045 ;
        RECT 110.080 46.000 110.220 47.500 ;
        RECT 120.685 47.360 120.975 47.405 ;
        RECT 123.805 47.360 124.095 47.405 ;
        RECT 125.695 47.360 125.985 47.405 ;
        RECT 129.310 47.360 129.630 47.420 ;
        RECT 120.685 47.220 125.985 47.360 ;
        RECT 120.685 47.175 120.975 47.220 ;
        RECT 123.805 47.175 124.095 47.220 ;
        RECT 125.695 47.175 125.985 47.220 ;
        RECT 126.180 47.220 129.630 47.360 ;
        RECT 125.185 47.020 125.475 47.065 ;
        RECT 126.180 47.020 126.320 47.220 ;
        RECT 129.310 47.160 129.630 47.220 ;
        RECT 125.185 46.880 126.320 47.020 ;
        RECT 126.565 47.020 126.855 47.065 ;
        RECT 130.690 47.020 131.010 47.080 ;
        RECT 126.565 46.880 131.010 47.020 ;
        RECT 125.185 46.835 125.475 46.880 ;
        RECT 126.565 46.835 126.855 46.880 ;
        RECT 130.690 46.820 131.010 46.880 ;
        RECT 119.605 46.385 119.895 46.700 ;
        RECT 120.685 46.680 120.975 46.725 ;
        RECT 124.265 46.680 124.555 46.725 ;
        RECT 126.100 46.680 126.390 46.725 ;
        RECT 127.025 46.680 127.315 46.725 ;
        RECT 120.685 46.540 126.390 46.680 ;
        RECT 120.685 46.495 120.975 46.540 ;
        RECT 124.265 46.495 124.555 46.540 ;
        RECT 126.100 46.495 126.390 46.540 ;
        RECT 126.640 46.540 127.315 46.680 ;
        RECT 126.640 46.400 126.780 46.540 ;
        RECT 127.025 46.495 127.315 46.540 ;
        RECT 117.365 46.340 117.655 46.385 ;
        RECT 119.305 46.340 119.895 46.385 ;
        RECT 122.545 46.340 123.195 46.385 ;
        RECT 117.365 46.200 118.960 46.340 ;
        RECT 117.365 46.155 117.655 46.200 ;
        RECT 108.165 45.860 110.220 46.000 ;
        RECT 118.820 46.000 118.960 46.200 ;
        RECT 119.305 46.200 123.560 46.340 ;
        RECT 119.305 46.155 119.595 46.200 ;
        RECT 122.545 46.155 123.195 46.200 ;
        RECT 120.570 46.000 120.890 46.060 ;
        RECT 118.820 45.860 120.890 46.000 ;
        RECT 123.420 46.000 123.560 46.200 ;
        RECT 126.550 46.140 126.870 46.400 ;
        RECT 127.485 46.155 127.775 46.385 ;
        RECT 127.560 46.000 127.700 46.155 ;
        RECT 123.420 45.860 127.700 46.000 ;
        RECT 108.165 45.815 108.455 45.860 ;
        RECT 120.570 45.800 120.890 45.860 ;
        RECT 88.980 45.180 152.240 45.660 ;
        RECT 88.980 40.220 89.460 45.180 ;
        RECT 99.425 44.980 99.715 45.025 ;
        RECT 100.790 44.980 101.110 45.040 ;
        RECT 99.425 44.840 101.110 44.980 ;
        RECT 99.425 44.795 99.715 44.840 ;
        RECT 100.790 44.780 101.110 44.840 ;
        RECT 110.450 44.780 110.770 45.040 ;
        RECT 111.830 44.980 112.150 45.040 ;
        RECT 112.305 44.980 112.595 45.025 ;
        RECT 111.830 44.840 112.595 44.980 ;
        RECT 111.830 44.780 112.150 44.840 ;
        RECT 112.305 44.795 112.595 44.840 ;
        RECT 114.145 44.980 114.435 45.025 ;
        RECT 115.050 44.980 115.370 45.040 ;
        RECT 114.145 44.840 115.370 44.980 ;
        RECT 114.145 44.795 114.435 44.840 ;
        RECT 115.050 44.780 115.370 44.840 ;
        RECT 129.310 44.780 129.630 45.040 ;
        RECT 131.150 44.780 131.470 45.040 ;
        RECT 134.370 44.780 134.690 45.040 ;
        RECT 134.830 44.780 135.150 45.040 ;
        RECT 137.605 44.980 137.895 45.025 ;
        RECT 137.605 44.840 140.580 44.980 ;
        RECT 137.605 44.795 137.895 44.840 ;
        RECT 97.110 44.640 97.430 44.700 ;
        RECT 97.585 44.640 97.875 44.685 ;
        RECT 97.110 44.500 97.875 44.640 ;
        RECT 97.110 44.440 97.430 44.500 ;
        RECT 97.585 44.455 97.875 44.500 ;
        RECT 100.345 44.640 100.635 44.685 ;
        RECT 104.485 44.640 104.775 44.685 ;
        RECT 100.345 44.500 104.775 44.640 ;
        RECT 100.345 44.455 100.635 44.500 ;
        RECT 104.485 44.455 104.775 44.500 ;
        RECT 105.850 44.640 106.170 44.700 ;
        RECT 106.325 44.640 106.615 44.685 ;
        RECT 111.385 44.640 111.675 44.685 ;
        RECT 105.850 44.500 111.675 44.640 ;
        RECT 96.205 44.115 96.495 44.345 ;
        RECT 96.280 43.340 96.420 44.115 ;
        RECT 97.660 43.960 97.800 44.455 ;
        RECT 105.850 44.440 106.170 44.500 ;
        RECT 106.325 44.455 106.615 44.500 ;
        RECT 111.385 44.455 111.675 44.500 ;
        RECT 113.210 44.440 113.530 44.700 ;
        RECT 127.010 44.685 127.330 44.700 ;
        RECT 126.895 44.455 127.330 44.685 ;
        RECT 131.240 44.640 131.380 44.780 ;
        RECT 131.240 44.500 132.300 44.640 ;
        RECT 127.010 44.440 127.330 44.455 ;
        RECT 102.185 44.300 102.475 44.345 ;
        RECT 104.010 44.300 104.330 44.360 ;
        RECT 102.185 44.160 104.330 44.300 ;
        RECT 102.185 44.115 102.475 44.160 ;
        RECT 104.010 44.100 104.330 44.160 ;
        RECT 105.390 44.300 105.710 44.360 ;
        RECT 111.845 44.300 112.135 44.345 ;
        RECT 105.390 44.160 112.135 44.300 ;
        RECT 105.390 44.100 105.710 44.160 ;
        RECT 111.845 44.115 112.135 44.160 ;
        RECT 114.605 44.115 114.895 44.345 ;
        RECT 120.110 44.300 120.430 44.360 ;
        RECT 122.425 44.300 122.715 44.345 ;
        RECT 120.110 44.160 122.715 44.300 ;
        RECT 114.680 43.960 114.820 44.115 ;
        RECT 120.110 44.100 120.430 44.160 ;
        RECT 122.425 44.115 122.715 44.160 ;
        RECT 127.485 44.115 127.775 44.345 ;
        RECT 97.660 43.820 114.820 43.960 ;
        RECT 125.645 43.960 125.935 44.005 ;
        RECT 126.105 43.960 126.395 44.005 ;
        RECT 125.645 43.820 126.395 43.960 ;
        RECT 125.645 43.775 125.935 43.820 ;
        RECT 126.105 43.775 126.395 43.820 ;
        RECT 127.010 43.960 127.330 44.020 ;
        RECT 127.560 43.960 127.700 44.115 ;
        RECT 127.930 44.100 128.250 44.360 ;
        RECT 128.405 44.300 128.695 44.345 ;
        RECT 131.610 44.300 131.930 44.360 ;
        RECT 132.160 44.345 132.300 44.500 ;
        RECT 134.460 44.345 134.600 44.780 ;
        RECT 128.405 44.160 131.930 44.300 ;
        RECT 128.405 44.115 128.695 44.160 ;
        RECT 131.610 44.100 131.930 44.160 ;
        RECT 132.085 44.115 132.375 44.345 ;
        RECT 134.385 44.115 134.675 44.345 ;
        RECT 134.920 44.300 135.060 44.780 ;
        RECT 138.065 44.640 138.355 44.685 ;
        RECT 136.760 44.500 138.355 44.640 ;
        RECT 136.760 44.345 136.900 44.500 ;
        RECT 138.065 44.455 138.355 44.500 ;
        RECT 138.970 44.440 139.290 44.700 ;
        RECT 140.440 44.685 140.580 44.840 ;
        RECT 142.205 44.795 142.495 45.025 ;
        RECT 140.365 44.455 140.655 44.685 ;
        RECT 140.810 44.640 141.130 44.700 ;
        RECT 141.365 44.640 141.655 44.685 ;
        RECT 140.810 44.500 141.655 44.640 ;
        RECT 136.685 44.300 136.975 44.345 ;
        RECT 134.920 44.160 136.975 44.300 ;
        RECT 136.685 44.115 136.975 44.160 ;
        RECT 137.605 44.300 137.895 44.345 ;
        RECT 139.060 44.300 139.200 44.440 ;
        RECT 137.605 44.160 139.200 44.300 ;
        RECT 140.440 44.300 140.580 44.455 ;
        RECT 140.810 44.440 141.130 44.500 ;
        RECT 141.365 44.455 141.655 44.500 ;
        RECT 142.280 44.300 142.420 44.795 ;
        RECT 144.045 44.300 144.335 44.345 ;
        RECT 140.440 44.160 141.960 44.300 ;
        RECT 142.280 44.160 144.335 44.300 ;
        RECT 137.605 44.115 137.895 44.160 ;
        RECT 134.830 43.960 135.150 44.020 ;
        RECT 127.010 43.820 135.150 43.960 ;
        RECT 127.010 43.760 127.330 43.820 ;
        RECT 134.830 43.760 135.150 43.820 ;
        RECT 141.820 43.340 141.960 44.160 ;
        RECT 144.045 44.115 144.335 44.160 ;
        RECT 146.345 44.115 146.635 44.345 ;
        RECT 142.650 43.960 142.970 44.020 ;
        RECT 146.420 43.960 146.560 44.115 ;
        RECT 142.650 43.820 146.560 43.960 ;
        RECT 142.650 43.760 142.970 43.820 ;
        RECT 96.190 43.080 96.510 43.340 ;
        RECT 100.345 43.280 100.635 43.325 ;
        RECT 107.230 43.280 107.550 43.340 ;
        RECT 100.345 43.140 107.550 43.280 ;
        RECT 100.345 43.095 100.635 43.140 ;
        RECT 107.230 43.080 107.550 43.140 ;
        RECT 126.550 43.280 126.870 43.340 ;
        RECT 131.625 43.280 131.915 43.325 ;
        RECT 126.550 43.140 131.915 43.280 ;
        RECT 126.550 43.080 126.870 43.140 ;
        RECT 131.625 43.095 131.915 43.140 ;
        RECT 133.925 43.280 134.215 43.325 ;
        RECT 134.370 43.280 134.690 43.340 ;
        RECT 133.925 43.140 134.690 43.280 ;
        RECT 133.925 43.095 134.215 43.140 ;
        RECT 134.370 43.080 134.690 43.140 ;
        RECT 139.905 43.280 140.195 43.325 ;
        RECT 141.285 43.280 141.575 43.325 ;
        RECT 139.905 43.140 141.575 43.280 ;
        RECT 139.905 43.095 140.195 43.140 ;
        RECT 141.285 43.095 141.575 43.140 ;
        RECT 141.730 43.080 142.050 43.340 ;
        RECT 143.110 43.080 143.430 43.340 ;
        RECT 146.330 43.280 146.650 43.340 ;
        RECT 146.805 43.280 147.095 43.325 ;
        RECT 146.330 43.140 147.095 43.280 ;
        RECT 146.330 43.080 146.650 43.140 ;
        RECT 146.805 43.095 147.095 43.140 ;
        RECT 152.900 42.940 153.380 47.900 ;
        RECT 91.060 42.460 153.380 42.940 ;
        RECT 131.610 42.260 131.930 42.320 ;
        RECT 138.985 42.260 139.275 42.305 ;
        RECT 142.650 42.260 142.970 42.320 ;
        RECT 149.550 42.260 149.870 42.320 ;
        RECT 131.610 42.120 139.275 42.260 ;
        RECT 131.610 42.060 131.930 42.120 ;
        RECT 138.985 42.075 139.275 42.120 ;
        RECT 141.820 42.120 149.870 42.260 ;
        RECT 141.820 41.920 141.960 42.120 ;
        RECT 142.650 42.060 142.970 42.120 ;
        RECT 149.550 42.060 149.870 42.120 ;
        RECT 109.620 41.780 141.960 41.920 ;
        RECT 142.155 41.920 142.445 41.965 ;
        RECT 144.045 41.920 144.335 41.965 ;
        RECT 147.165 41.920 147.455 41.965 ;
        RECT 142.155 41.780 147.455 41.920 ;
        RECT 109.620 41.640 109.760 41.780 ;
        RECT 142.155 41.735 142.445 41.780 ;
        RECT 144.045 41.735 144.335 41.780 ;
        RECT 147.165 41.735 147.455 41.780 ;
        RECT 100.345 41.580 100.635 41.625 ;
        RECT 109.530 41.580 109.850 41.640 ;
        RECT 100.345 41.440 109.850 41.580 ;
        RECT 100.345 41.395 100.635 41.440 ;
        RECT 109.530 41.380 109.850 41.440 ;
        RECT 142.665 41.580 142.955 41.625 ;
        RECT 143.110 41.580 143.430 41.640 ;
        RECT 142.665 41.440 143.430 41.580 ;
        RECT 142.665 41.395 142.955 41.440 ;
        RECT 143.110 41.380 143.430 41.440 ;
        RECT 90.210 41.240 90.530 41.300 ;
        RECT 92.525 41.240 92.815 41.285 ;
        RECT 90.210 41.100 92.815 41.240 ;
        RECT 90.210 41.040 90.530 41.100 ;
        RECT 92.525 41.055 92.815 41.100 ;
        RECT 98.965 41.055 99.255 41.285 ;
        RECT 93.445 40.560 93.735 40.605 ;
        RECT 96.190 40.560 96.510 40.620 ;
        RECT 99.040 40.560 99.180 41.055 ;
        RECT 138.970 41.040 139.290 41.300 ;
        RECT 139.905 41.240 140.195 41.285 ;
        RECT 139.905 41.100 141.040 41.240 ;
        RECT 139.905 41.055 140.195 41.100 ;
        RECT 139.060 40.900 139.200 41.040 ;
        RECT 140.350 40.900 140.670 40.960 ;
        RECT 139.060 40.760 140.670 40.900 ;
        RECT 140.350 40.700 140.670 40.760 ;
        RECT 140.900 40.620 141.040 41.100 ;
        RECT 141.270 41.040 141.590 41.300 ;
        RECT 141.750 41.240 142.040 41.285 ;
        RECT 143.585 41.240 143.875 41.285 ;
        RECT 147.165 41.240 147.455 41.285 ;
        RECT 141.750 41.100 147.455 41.240 ;
        RECT 141.750 41.055 142.040 41.100 ;
        RECT 143.585 41.055 143.875 41.100 ;
        RECT 147.165 41.055 147.455 41.100 ;
        RECT 144.945 40.900 145.595 40.945 ;
        RECT 146.330 40.900 146.650 40.960 ;
        RECT 148.245 40.945 148.535 41.260 ;
        RECT 148.245 40.900 148.835 40.945 ;
        RECT 144.945 40.760 148.835 40.900 ;
        RECT 144.945 40.715 145.595 40.760 ;
        RECT 146.330 40.700 146.650 40.760 ;
        RECT 148.545 40.715 148.835 40.760 ;
        RECT 93.445 40.420 99.180 40.560 ;
        RECT 93.445 40.375 93.735 40.420 ;
        RECT 96.190 40.360 96.510 40.420 ;
        RECT 140.810 40.360 141.130 40.620 ;
        RECT 142.190 40.560 142.510 40.620 ;
        RECT 150.025 40.560 150.315 40.605 ;
        RECT 142.190 40.420 150.315 40.560 ;
        RECT 142.190 40.360 142.510 40.420 ;
        RECT 150.025 40.375 150.315 40.420 ;
        RECT 88.980 39.740 152.240 40.220 ;
        RECT 0.995 35.915 2.505 36.290 ;
        RECT 0.995 35.560 59.410 35.915 ;
        RECT 0.995 35.135 2.505 35.560 ;
        RECT 59.055 34.420 59.410 35.560 ;
        RECT 88.980 34.780 89.460 39.740 ;
        RECT 99.500 39.400 101.480 39.540 ;
        RECT 99.500 38.860 99.640 39.400 ;
        RECT 95.820 38.720 99.640 38.860 ;
        RECT 95.820 38.580 95.960 38.720 ;
        RECT 99.885 38.675 100.175 38.905 ;
        RECT 101.340 38.860 101.480 39.400 ;
        RECT 102.170 39.340 102.490 39.600 ;
        RECT 106.310 39.340 106.630 39.600 ;
        RECT 107.780 39.400 116.660 39.540 ;
        RECT 107.230 38.860 107.550 38.920 ;
        RECT 101.340 38.720 107.550 38.860 ;
        RECT 95.730 38.320 96.050 38.580 ;
        RECT 96.650 38.520 96.970 38.580 ;
        RECT 98.950 38.520 99.270 38.580 ;
        RECT 96.650 38.380 99.270 38.520 ;
        RECT 99.960 38.520 100.100 38.675 ;
        RECT 107.230 38.660 107.550 38.720 ;
        RECT 104.010 38.520 104.330 38.580 ;
        RECT 107.780 38.520 107.920 39.400 ;
        RECT 113.685 39.200 113.975 39.245 ;
        RECT 115.510 39.200 115.830 39.260 ;
        RECT 113.685 39.060 115.830 39.200 ;
        RECT 113.685 39.015 113.975 39.060 ;
        RECT 115.510 39.000 115.830 39.060 ;
        RECT 108.165 38.860 108.455 38.905 ;
        RECT 108.165 38.720 108.840 38.860 ;
        RECT 108.165 38.675 108.455 38.720 ;
        RECT 99.960 38.380 104.330 38.520 ;
        RECT 96.650 38.320 96.970 38.380 ;
        RECT 98.950 38.320 99.270 38.380 ;
        RECT 104.010 38.320 104.330 38.380 ;
        RECT 104.560 38.380 107.920 38.520 ;
        RECT 108.700 38.520 108.840 38.720 ;
        RECT 109.530 38.660 109.850 38.920 ;
        RECT 109.990 38.660 110.310 38.920 ;
        RECT 110.925 38.860 111.215 38.905 ;
        RECT 114.145 38.860 114.435 38.905 ;
        RECT 110.925 38.720 114.435 38.860 ;
        RECT 116.520 38.860 116.660 39.400 ;
        RECT 121.490 39.340 121.810 39.600 ;
        RECT 121.950 39.340 122.270 39.600 ;
        RECT 136.685 39.540 136.975 39.585 ;
        RECT 139.890 39.540 140.210 39.600 ;
        RECT 123.880 39.400 130.920 39.540 ;
        RECT 121.580 38.905 121.720 39.340 ;
        RECT 122.040 39.200 122.180 39.340 ;
        RECT 123.880 39.245 124.020 39.400 ;
        RECT 123.805 39.200 124.095 39.245 ;
        RECT 122.040 39.060 124.095 39.200 ;
        RECT 123.805 39.015 124.095 39.060 ;
        RECT 125.260 39.060 128.160 39.200 ;
        RECT 120.125 38.860 120.415 38.905 ;
        RECT 116.520 38.720 120.415 38.860 ;
        RECT 110.925 38.675 111.215 38.720 ;
        RECT 114.145 38.675 114.435 38.720 ;
        RECT 120.125 38.675 120.415 38.720 ;
        RECT 121.505 38.675 121.795 38.905 ;
        RECT 122.410 38.660 122.730 38.920 ;
        RECT 123.330 38.660 123.650 38.920 ;
        RECT 124.250 38.660 124.570 38.920 ;
        RECT 112.290 38.520 112.610 38.580 ;
        RECT 108.700 38.380 112.610 38.520 ;
        RECT 98.505 38.180 98.795 38.225 ;
        RECT 100.790 38.180 101.110 38.240 ;
        RECT 98.505 38.040 101.110 38.180 ;
        RECT 98.505 37.995 98.795 38.040 ;
        RECT 100.790 37.980 101.110 38.040 ;
        RECT 103.550 38.180 103.870 38.240 ;
        RECT 104.560 38.180 104.700 38.380 ;
        RECT 103.550 38.040 104.700 38.180 ;
        RECT 105.390 38.180 105.710 38.240 ;
        RECT 105.865 38.180 106.155 38.225 ;
        RECT 108.700 38.180 108.840 38.380 ;
        RECT 112.290 38.320 112.610 38.380 ;
        RECT 114.605 38.520 114.895 38.565 ;
        RECT 115.050 38.520 115.370 38.580 ;
        RECT 114.605 38.380 115.370 38.520 ;
        RECT 114.605 38.335 114.895 38.380 ;
        RECT 115.050 38.320 115.370 38.380 ;
        RECT 115.525 38.520 115.815 38.565 ;
        RECT 115.970 38.520 116.290 38.580 ;
        RECT 115.525 38.380 116.290 38.520 ;
        RECT 115.525 38.335 115.815 38.380 ;
        RECT 115.970 38.320 116.290 38.380 ;
        RECT 117.810 38.520 118.130 38.580 ;
        RECT 119.205 38.520 119.495 38.565 ;
        RECT 117.810 38.380 119.495 38.520 ;
        RECT 117.810 38.320 118.130 38.380 ;
        RECT 119.205 38.335 119.495 38.380 ;
        RECT 119.650 38.520 119.970 38.580 ;
        RECT 125.260 38.520 125.400 39.060 ;
        RECT 125.630 38.660 125.950 38.920 ;
        RECT 126.090 38.860 126.410 38.920 ;
        RECT 126.565 38.860 126.855 38.905 ;
        RECT 126.090 38.720 126.855 38.860 ;
        RECT 126.090 38.660 126.410 38.720 ;
        RECT 126.565 38.675 126.855 38.720 ;
        RECT 127.025 38.675 127.315 38.905 ;
        RECT 119.650 38.380 125.400 38.520 ;
        RECT 127.100 38.520 127.240 38.675 ;
        RECT 127.470 38.660 127.790 38.920 ;
        RECT 128.020 38.860 128.160 39.060 ;
        RECT 129.400 39.060 130.460 39.200 ;
        RECT 128.865 38.860 129.155 38.905 ;
        RECT 128.020 38.720 129.155 38.860 ;
        RECT 128.865 38.675 129.155 38.720 ;
        RECT 129.400 38.520 129.540 39.060 ;
        RECT 129.785 38.675 130.075 38.905 ;
        RECT 127.100 38.380 129.540 38.520 ;
        RECT 119.650 38.320 119.970 38.380 ;
        RECT 105.390 38.040 108.840 38.180 ;
        RECT 103.550 37.980 103.870 38.040 ;
        RECT 105.390 37.980 105.710 38.040 ;
        RECT 105.865 37.995 106.155 38.040 ;
        RECT 111.830 37.980 112.150 38.240 ;
        RECT 112.750 38.180 113.070 38.240 ;
        RECT 120.585 38.180 120.875 38.225 ;
        RECT 112.750 38.040 120.875 38.180 ;
        RECT 112.750 37.980 113.070 38.040 ;
        RECT 120.585 37.995 120.875 38.040 ;
        RECT 121.030 37.980 121.350 38.240 ;
        RECT 121.490 38.180 121.810 38.240 ;
        RECT 125.185 38.180 125.475 38.225 ;
        RECT 129.860 38.180 130.000 38.675 ;
        RECT 130.320 38.520 130.460 39.060 ;
        RECT 130.780 38.860 130.920 39.400 ;
        RECT 136.685 39.400 140.210 39.540 ;
        RECT 136.685 39.355 136.975 39.400 ;
        RECT 139.890 39.340 140.210 39.400 ;
        RECT 140.350 39.540 140.670 39.600 ;
        RECT 142.190 39.540 142.510 39.600 ;
        RECT 140.350 39.400 142.510 39.540 ;
        RECT 140.350 39.340 140.670 39.400 ;
        RECT 142.190 39.340 142.510 39.400 ;
        RECT 140.810 39.200 141.130 39.260 ;
        RECT 141.285 39.200 141.575 39.245 ;
        RECT 140.810 39.060 150.240 39.200 ;
        RECT 140.810 39.000 141.130 39.060 ;
        RECT 141.285 39.015 141.575 39.060 ;
        RECT 150.100 38.920 150.240 39.060 ;
        RECT 132.545 38.860 132.835 38.905 ;
        RECT 130.780 38.720 132.835 38.860 ;
        RECT 132.545 38.675 132.835 38.720 ;
        RECT 134.370 38.660 134.690 38.920 ;
        RECT 134.830 38.860 135.150 38.920 ;
        RECT 137.435 38.860 137.725 38.905 ;
        RECT 134.830 38.720 137.820 38.860 ;
        RECT 134.830 38.660 135.150 38.720 ;
        RECT 137.435 38.675 137.820 38.720 ;
        RECT 134.460 38.520 134.600 38.660 ;
        RECT 130.320 38.380 134.600 38.520 ;
        RECT 137.680 38.240 137.820 38.675 ;
        RECT 139.890 38.660 140.210 38.920 ;
        RECT 144.045 38.860 144.335 38.905 ;
        RECT 147.265 38.860 147.555 38.905 ;
        RECT 144.045 38.720 147.555 38.860 ;
        RECT 144.045 38.675 144.335 38.720 ;
        RECT 147.265 38.675 147.555 38.720 ;
        RECT 150.010 38.660 150.330 38.920 ;
        RECT 138.970 38.320 139.290 38.580 ;
        RECT 139.445 38.335 139.735 38.565 ;
        RECT 141.730 38.520 142.050 38.580 ;
        RECT 143.585 38.520 143.875 38.565 ;
        RECT 141.730 38.380 143.875 38.520 ;
        RECT 121.490 38.040 124.940 38.180 ;
        RECT 121.490 37.980 121.810 38.040 ;
        RECT 98.965 37.840 99.255 37.885 ;
        RECT 99.870 37.840 100.190 37.900 ;
        RECT 98.965 37.700 100.190 37.840 ;
        RECT 98.965 37.655 99.255 37.700 ;
        RECT 99.870 37.640 100.190 37.700 ;
        RECT 101.265 37.840 101.555 37.885 ;
        RECT 104.930 37.840 105.250 37.900 ;
        RECT 101.265 37.700 105.250 37.840 ;
        RECT 101.265 37.655 101.555 37.700 ;
        RECT 104.930 37.640 105.250 37.700 ;
        RECT 108.625 37.840 108.915 37.885 ;
        RECT 110.910 37.840 111.230 37.900 ;
        RECT 108.625 37.700 111.230 37.840 ;
        RECT 108.625 37.655 108.915 37.700 ;
        RECT 110.910 37.640 111.230 37.700 ;
        RECT 111.370 37.640 111.690 37.900 ;
        RECT 115.065 37.840 115.355 37.885 ;
        RECT 118.730 37.840 119.050 37.900 ;
        RECT 115.065 37.700 119.050 37.840 ;
        RECT 115.065 37.655 115.355 37.700 ;
        RECT 118.730 37.640 119.050 37.700 ;
        RECT 120.110 37.840 120.430 37.900 ;
        RECT 123.330 37.840 123.650 37.900 ;
        RECT 120.110 37.700 123.650 37.840 ;
        RECT 124.800 37.840 124.940 38.040 ;
        RECT 125.185 38.040 130.000 38.180 ;
        RECT 125.185 37.995 125.475 38.040 ;
        RECT 131.150 37.980 131.470 38.240 ;
        RECT 131.610 38.180 131.930 38.240 ;
        RECT 131.610 38.040 137.360 38.180 ;
        RECT 131.610 37.980 131.930 38.040 ;
        RECT 127.470 37.840 127.790 37.900 ;
        RECT 124.800 37.700 127.790 37.840 ;
        RECT 120.110 37.640 120.430 37.700 ;
        RECT 123.330 37.640 123.650 37.700 ;
        RECT 127.470 37.640 127.790 37.700 ;
        RECT 127.930 37.840 128.250 37.900 ;
        RECT 128.405 37.840 128.695 37.885 ;
        RECT 127.930 37.700 128.695 37.840 ;
        RECT 127.930 37.640 128.250 37.700 ;
        RECT 128.405 37.655 128.695 37.700 ;
        RECT 129.785 37.840 130.075 37.885 ;
        RECT 130.230 37.840 130.550 37.900 ;
        RECT 129.785 37.700 130.550 37.840 ;
        RECT 129.785 37.655 130.075 37.700 ;
        RECT 130.230 37.640 130.550 37.700 ;
        RECT 130.690 37.840 131.010 37.900 ;
        RECT 132.085 37.840 132.375 37.885 ;
        RECT 130.690 37.700 132.375 37.840 ;
        RECT 137.220 37.840 137.360 38.040 ;
        RECT 137.590 37.980 137.910 38.240 ;
        RECT 139.520 38.180 139.660 38.335 ;
        RECT 141.730 38.320 142.050 38.380 ;
        RECT 143.585 38.335 143.875 38.380 ;
        RECT 141.285 38.180 141.575 38.225 ;
        RECT 139.520 38.040 141.575 38.180 ;
        RECT 141.285 37.995 141.575 38.040 ;
        RECT 139.430 37.840 139.750 37.900 ;
        RECT 137.220 37.700 139.750 37.840 ;
        RECT 130.690 37.640 131.010 37.700 ;
        RECT 132.085 37.655 132.375 37.700 ;
        RECT 139.430 37.640 139.750 37.700 ;
        RECT 145.870 37.640 146.190 37.900 ;
        RECT 152.900 37.500 153.380 42.460 ;
        RECT 91.060 37.020 153.380 37.500 ;
        RECT 93.905 36.820 94.195 36.865 ;
        RECT 97.125 36.820 97.415 36.865 ;
        RECT 93.905 36.680 97.415 36.820 ;
        RECT 93.905 36.635 94.195 36.680 ;
        RECT 97.125 36.635 97.415 36.680 ;
        RECT 98.965 36.820 99.255 36.865 ;
        RECT 99.870 36.820 100.190 36.880 ;
        RECT 108.165 36.820 108.455 36.865 ;
        RECT 109.530 36.820 109.850 36.880 ;
        RECT 98.965 36.680 106.540 36.820 ;
        RECT 98.965 36.635 99.255 36.680 ;
        RECT 95.285 36.480 95.575 36.525 ;
        RECT 96.650 36.480 96.970 36.540 ;
        RECT 95.285 36.340 96.970 36.480 ;
        RECT 95.285 36.295 95.575 36.340 ;
        RECT 92.525 35.800 92.815 35.845 ;
        RECT 93.430 35.800 93.750 35.860 ;
        RECT 95.360 35.800 95.500 36.295 ;
        RECT 96.650 36.280 96.970 36.340 ;
        RECT 95.730 35.940 96.050 36.200 ;
        RECT 97.200 36.140 97.340 36.635 ;
        RECT 99.870 36.620 100.190 36.680 ;
        RECT 98.045 36.480 98.335 36.525 ;
        RECT 98.045 36.340 101.940 36.480 ;
        RECT 98.045 36.295 98.335 36.340 ;
        RECT 100.330 36.140 100.650 36.200 ;
        RECT 97.200 36.000 100.650 36.140 ;
        RECT 100.330 35.940 100.650 36.000 ;
        RECT 92.525 35.660 95.500 35.800 ;
        RECT 95.820 35.800 95.960 35.940 ;
        RECT 98.505 35.800 98.795 35.845 ;
        RECT 95.820 35.660 98.795 35.800 ;
        RECT 92.525 35.615 92.815 35.660 ;
        RECT 93.430 35.600 93.750 35.660 ;
        RECT 98.505 35.615 98.795 35.660 ;
        RECT 100.790 35.600 101.110 35.860 ;
        RECT 100.345 35.460 100.635 35.505 ;
        RECT 94.900 35.320 100.635 35.460 ;
        RECT 101.800 35.460 101.940 36.340 ;
        RECT 102.170 36.280 102.490 36.540 ;
        RECT 103.105 36.480 103.395 36.525 ;
        RECT 103.105 36.340 106.080 36.480 ;
        RECT 103.105 36.295 103.395 36.340 ;
        RECT 102.260 36.140 102.400 36.280 ;
        RECT 105.940 36.200 106.080 36.340 ;
        RECT 102.260 36.000 104.700 36.140 ;
        RECT 102.645 35.800 102.935 35.845 ;
        RECT 103.550 35.800 103.870 35.860 ;
        RECT 104.560 35.845 104.700 36.000 ;
        RECT 105.850 35.940 106.170 36.200 ;
        RECT 106.400 36.185 106.540 36.680 ;
        RECT 108.165 36.680 109.850 36.820 ;
        RECT 108.165 36.635 108.455 36.680 ;
        RECT 109.530 36.620 109.850 36.680 ;
        RECT 110.910 36.620 111.230 36.880 ;
        RECT 113.225 36.820 113.515 36.865 ;
        RECT 119.650 36.820 119.970 36.880 ;
        RECT 113.225 36.680 119.970 36.820 ;
        RECT 113.225 36.635 113.515 36.680 ;
        RECT 119.650 36.620 119.970 36.680 ;
        RECT 120.585 36.635 120.875 36.865 ;
        RECT 121.030 36.820 121.350 36.880 ;
        RECT 122.425 36.820 122.715 36.865 ;
        RECT 121.030 36.680 122.715 36.820 ;
        RECT 106.325 35.955 106.615 36.185 ;
        RECT 111.000 36.140 111.140 36.620 ;
        RECT 115.065 36.480 115.355 36.525 ;
        RECT 115.970 36.480 116.290 36.540 ;
        RECT 120.110 36.480 120.430 36.540 ;
        RECT 115.065 36.340 116.290 36.480 ;
        RECT 115.065 36.295 115.355 36.340 ;
        RECT 115.970 36.280 116.290 36.340 ;
        RECT 116.980 36.340 120.430 36.480 ;
        RECT 120.660 36.480 120.800 36.635 ;
        RECT 121.030 36.620 121.350 36.680 ;
        RECT 122.425 36.635 122.715 36.680 ;
        RECT 125.630 36.820 125.950 36.880 ;
        RECT 130.245 36.820 130.535 36.865 ;
        RECT 131.610 36.820 131.930 36.880 ;
        RECT 136.685 36.820 136.975 36.865 ;
        RECT 138.970 36.820 139.290 36.880 ;
        RECT 125.630 36.680 130.535 36.820 ;
        RECT 125.630 36.620 125.950 36.680 ;
        RECT 130.245 36.635 130.535 36.680 ;
        RECT 131.240 36.680 131.930 36.820 ;
        RECT 120.660 36.340 128.620 36.480 ;
        RECT 111.385 36.140 111.675 36.185 ;
        RECT 112.750 36.140 113.070 36.200 ;
        RECT 114.145 36.140 114.435 36.185 ;
        RECT 111.000 36.000 114.435 36.140 ;
        RECT 111.385 35.955 111.675 36.000 ;
        RECT 112.750 35.940 113.070 36.000 ;
        RECT 114.145 35.955 114.435 36.000 ;
        RECT 115.510 35.940 115.830 36.200 ;
        RECT 116.980 36.140 117.120 36.340 ;
        RECT 120.110 36.280 120.430 36.340 ;
        RECT 116.060 36.000 117.120 36.140 ;
        RECT 117.365 36.140 117.655 36.185 ;
        RECT 117.365 36.000 120.340 36.140 ;
        RECT 102.645 35.660 103.870 35.800 ;
        RECT 102.645 35.615 102.935 35.660 ;
        RECT 103.550 35.600 103.870 35.660 ;
        RECT 104.485 35.615 104.775 35.845 ;
        RECT 105.405 35.615 105.695 35.845 ;
        RECT 105.480 35.460 105.620 35.615 ;
        RECT 107.230 35.600 107.550 35.860 ;
        RECT 109.530 35.600 109.850 35.860 ;
        RECT 110.465 35.615 110.755 35.845 ;
        RECT 101.800 35.320 105.620 35.460 ;
        RECT 94.900 35.165 95.040 35.320 ;
        RECT 100.345 35.275 100.635 35.320 ;
        RECT 94.825 34.935 95.115 35.165 ;
        RECT 95.730 35.120 96.050 35.180 ;
        RECT 97.125 35.120 97.415 35.165 ;
        RECT 95.730 34.980 97.415 35.120 ;
        RECT 95.730 34.920 96.050 34.980 ;
        RECT 97.125 34.935 97.415 34.980 ;
        RECT 99.870 34.920 100.190 35.180 ;
        RECT 102.185 35.120 102.475 35.165 ;
        RECT 110.540 35.120 110.680 35.615 ;
        RECT 110.910 35.600 111.230 35.860 ;
        RECT 111.830 35.800 112.150 35.860 ;
        RECT 112.305 35.800 112.595 35.845 ;
        RECT 111.830 35.660 112.595 35.800 ;
        RECT 111.830 35.600 112.150 35.660 ;
        RECT 112.305 35.615 112.595 35.660 ;
        RECT 114.605 35.800 114.895 35.845 ;
        RECT 115.600 35.800 115.740 35.940 ;
        RECT 116.060 35.860 116.200 36.000 ;
        RECT 117.365 35.955 117.655 36.000 ;
        RECT 114.605 35.660 115.740 35.800 ;
        RECT 114.605 35.615 114.895 35.660 ;
        RECT 112.380 35.460 112.520 35.615 ;
        RECT 115.970 35.600 116.290 35.860 ;
        RECT 116.445 35.615 116.735 35.845 ;
        RECT 117.825 35.800 118.115 35.845 ;
        RECT 119.190 35.800 119.510 35.860 ;
        RECT 117.825 35.660 119.510 35.800 ;
        RECT 120.200 35.800 120.340 36.000 ;
        RECT 121.030 35.940 121.350 36.200 ;
        RECT 121.950 36.140 122.270 36.200 ;
        RECT 121.950 36.000 123.100 36.140 ;
        RECT 121.950 35.940 122.270 36.000 ;
        RECT 120.200 35.660 120.800 35.800 ;
        RECT 117.825 35.615 118.115 35.660 ;
        RECT 116.525 35.460 116.665 35.615 ;
        RECT 112.380 35.320 116.665 35.460 ;
        RECT 102.185 34.980 110.680 35.120 ;
        RECT 114.590 35.120 114.910 35.180 ;
        RECT 117.900 35.120 118.040 35.615 ;
        RECT 119.190 35.600 119.510 35.660 ;
        RECT 120.110 35.260 120.430 35.520 ;
        RECT 120.660 35.460 120.800 35.660 ;
        RECT 121.490 35.600 121.810 35.860 ;
        RECT 122.960 35.800 123.100 36.000 ;
        RECT 124.250 35.940 124.570 36.200 ;
        RECT 123.510 35.800 123.800 35.845 ;
        RECT 122.960 35.660 123.800 35.800 ;
        RECT 123.510 35.615 123.800 35.660 ;
        RECT 124.340 35.460 124.480 35.940 ;
        RECT 125.260 35.800 125.400 36.340 ;
        RECT 125.645 36.140 125.935 36.185 ;
        RECT 127.930 36.140 128.250 36.200 ;
        RECT 125.645 36.000 128.250 36.140 ;
        RECT 125.645 35.955 125.935 36.000 ;
        RECT 127.930 35.940 128.250 36.000 ;
        RECT 128.480 35.860 128.620 36.340 ;
        RECT 129.770 36.140 130.090 36.200 ;
        RECT 131.240 36.140 131.380 36.680 ;
        RECT 131.610 36.620 131.930 36.680 ;
        RECT 132.160 36.680 134.600 36.820 ;
        RECT 132.160 36.480 132.300 36.680 ;
        RECT 134.460 36.540 134.600 36.680 ;
        RECT 136.685 36.680 139.290 36.820 ;
        RECT 136.685 36.635 136.975 36.680 ;
        RECT 138.970 36.620 139.290 36.680 ;
        RECT 139.890 36.820 140.210 36.880 ;
        RECT 140.365 36.820 140.655 36.865 ;
        RECT 139.890 36.680 140.655 36.820 ;
        RECT 139.890 36.620 140.210 36.680 ;
        RECT 140.365 36.635 140.655 36.680 ;
        RECT 150.010 36.620 150.330 36.880 ;
        RECT 129.770 36.000 131.380 36.140 ;
        RECT 129.770 35.940 130.090 36.000 ;
        RECT 126.105 35.800 126.395 35.845 ;
        RECT 125.260 35.660 126.395 35.800 ;
        RECT 126.105 35.615 126.395 35.660 ;
        RECT 126.550 35.600 126.870 35.860 ;
        RECT 127.470 35.600 127.790 35.860 ;
        RECT 128.390 35.600 128.710 35.860 ;
        RECT 128.850 35.800 129.170 35.860 ;
        RECT 129.325 35.800 129.615 35.845 ;
        RECT 130.690 35.800 131.010 35.860 ;
        RECT 131.240 35.845 131.380 36.000 ;
        RECT 131.700 36.340 132.300 36.480 ;
        RECT 131.700 35.845 131.840 36.340 ;
        RECT 132.530 36.280 132.850 36.540 ;
        RECT 133.450 36.480 133.770 36.540 ;
        RECT 133.450 36.280 133.910 36.480 ;
        RECT 134.370 36.280 134.690 36.540 ;
        RECT 133.770 36.140 133.910 36.280 ;
        RECT 138.065 36.140 138.355 36.185 ;
        RECT 139.980 36.140 140.120 36.620 ;
        RECT 142.155 36.480 142.445 36.525 ;
        RECT 144.045 36.480 144.335 36.525 ;
        RECT 147.165 36.480 147.455 36.525 ;
        RECT 142.155 36.340 147.455 36.480 ;
        RECT 142.155 36.295 142.445 36.340 ;
        RECT 144.045 36.295 144.335 36.340 ;
        RECT 147.165 36.295 147.455 36.340 ;
        RECT 133.770 36.000 138.355 36.140 ;
        RECT 138.065 35.955 138.355 36.000 ;
        RECT 138.600 36.000 140.120 36.140 ;
        RECT 128.850 35.660 131.010 35.800 ;
        RECT 128.850 35.600 129.170 35.660 ;
        RECT 129.325 35.615 129.615 35.660 ;
        RECT 130.690 35.600 131.010 35.660 ;
        RECT 131.165 35.615 131.455 35.845 ;
        RECT 131.625 35.615 131.915 35.845 ;
        RECT 132.070 35.800 132.390 35.860 ;
        RECT 132.915 35.800 133.205 35.845 ;
        RECT 132.070 35.660 133.205 35.800 ;
        RECT 132.070 35.600 132.390 35.660 ;
        RECT 132.915 35.615 133.205 35.660 ;
        RECT 133.450 35.600 133.770 35.860 ;
        RECT 133.910 35.600 134.230 35.860 ;
        RECT 134.370 35.800 134.690 35.860 ;
        RECT 138.600 35.845 138.740 36.000 ;
        RECT 141.270 35.940 141.590 36.200 ;
        RECT 135.305 35.800 135.595 35.845 ;
        RECT 134.370 35.660 135.595 35.800 ;
        RECT 134.370 35.600 134.690 35.660 ;
        RECT 135.305 35.615 135.595 35.660 ;
        RECT 135.790 35.800 136.080 35.845 ;
        RECT 135.790 35.660 136.440 35.800 ;
        RECT 135.790 35.615 136.080 35.660 ;
        RECT 120.660 35.320 124.480 35.460 ;
        RECT 126.640 35.460 126.780 35.600 ;
        RECT 127.945 35.460 128.235 35.505 ;
        RECT 126.640 35.320 128.235 35.460 ;
        RECT 114.590 34.980 118.040 35.120 ;
        RECT 102.185 34.935 102.475 34.980 ;
        RECT 114.590 34.920 114.910 34.980 ;
        RECT 122.870 34.920 123.190 35.180 ;
        RECT 123.805 35.120 124.095 35.165 ;
        RECT 124.340 35.120 124.480 35.320 ;
        RECT 127.945 35.275 128.235 35.320 ;
        RECT 130.230 35.460 130.550 35.520 ;
        RECT 134.845 35.460 135.135 35.505 ;
        RECT 130.230 35.320 135.135 35.460 ;
        RECT 123.805 34.980 124.480 35.120 ;
        RECT 123.805 34.935 124.095 34.980 ;
        RECT 126.550 34.920 126.870 35.180 ;
        RECT 127.010 35.120 127.330 35.180 ;
        RECT 128.020 35.120 128.160 35.275 ;
        RECT 130.230 35.260 130.550 35.320 ;
        RECT 134.845 35.275 135.135 35.320 ;
        RECT 130.690 35.120 131.010 35.180 ;
        RECT 132.070 35.120 132.390 35.180 ;
        RECT 127.010 34.980 132.390 35.120 ;
        RECT 127.010 34.920 127.330 34.980 ;
        RECT 130.690 34.920 131.010 34.980 ;
        RECT 132.070 34.920 132.390 34.980 ;
        RECT 132.530 35.120 132.850 35.180 ;
        RECT 136.300 35.120 136.440 35.660 ;
        RECT 137.605 35.615 137.895 35.845 ;
        RECT 138.525 35.615 138.815 35.845 ;
        RECT 137.680 35.460 137.820 35.615 ;
        RECT 139.890 35.600 140.210 35.860 ;
        RECT 140.350 35.600 140.670 35.860 ;
        RECT 141.750 35.800 142.040 35.845 ;
        RECT 143.585 35.800 143.875 35.845 ;
        RECT 147.165 35.800 147.455 35.845 ;
        RECT 141.750 35.660 147.455 35.800 ;
        RECT 141.750 35.615 142.040 35.660 ;
        RECT 143.585 35.615 143.875 35.660 ;
        RECT 147.165 35.615 147.455 35.660 ;
        RECT 140.440 35.460 140.580 35.600 ;
        RECT 148.245 35.505 148.535 35.820 ;
        RECT 137.680 35.320 140.580 35.460 ;
        RECT 142.665 35.275 142.955 35.505 ;
        RECT 144.945 35.460 145.595 35.505 ;
        RECT 148.245 35.460 148.835 35.505 ;
        RECT 149.090 35.460 149.410 35.520 ;
        RECT 144.945 35.320 149.410 35.460 ;
        RECT 144.945 35.275 145.595 35.320 ;
        RECT 148.545 35.275 148.835 35.320 ;
        RECT 140.810 35.120 141.130 35.180 ;
        RECT 132.530 34.980 141.130 35.120 ;
        RECT 142.740 35.120 142.880 35.275 ;
        RECT 149.090 35.260 149.410 35.320 ;
        RECT 146.330 35.120 146.650 35.180 ;
        RECT 142.740 34.980 146.650 35.120 ;
        RECT 132.530 34.920 132.850 34.980 ;
        RECT 140.810 34.920 141.130 34.980 ;
        RECT 146.330 34.920 146.650 34.980 ;
        RECT 6.080 31.965 6.330 34.070 ;
        RECT 59.105 32.530 59.355 34.420 ;
        RECT 88.980 34.300 152.240 34.780 ;
        RECT 152.900 34.650 153.380 37.020 ;
        RECT 6.080 28.810 6.330 30.915 ;
        RECT 7.855 28.675 8.595 29.690 ;
        RECT 88.980 29.340 89.460 34.300 ;
        RECT 152.900 34.170 154.340 34.650 ;
        RECT 99.870 34.100 100.190 34.160 ;
        RECT 100.345 34.100 100.635 34.145 ;
        RECT 99.870 33.960 100.635 34.100 ;
        RECT 99.870 33.900 100.190 33.960 ;
        RECT 100.345 33.915 100.635 33.960 ;
        RECT 100.790 33.900 101.110 34.160 ;
        RECT 102.170 34.100 102.490 34.160 ;
        RECT 104.930 34.100 105.250 34.160 ;
        RECT 105.850 34.100 106.170 34.160 ;
        RECT 102.170 33.960 105.250 34.100 ;
        RECT 102.170 33.900 102.490 33.960 ;
        RECT 104.930 33.900 105.250 33.960 ;
        RECT 105.480 33.960 106.170 34.100 ;
        RECT 100.880 33.760 101.020 33.900 ;
        RECT 105.480 33.805 105.620 33.960 ;
        RECT 105.850 33.900 106.170 33.960 ;
        RECT 106.310 34.100 106.630 34.160 ;
        RECT 107.705 34.100 107.995 34.145 ;
        RECT 109.990 34.100 110.310 34.160 ;
        RECT 106.310 33.960 107.000 34.100 ;
        RECT 106.310 33.900 106.630 33.960 ;
        RECT 100.880 33.620 104.700 33.760 ;
        RECT 98.045 33.420 98.335 33.465 ;
        RECT 99.870 33.420 100.190 33.480 ;
        RECT 102.630 33.420 102.950 33.480 ;
        RECT 98.045 33.280 102.950 33.420 ;
        RECT 98.045 33.235 98.335 33.280 ;
        RECT 99.870 33.220 100.190 33.280 ;
        RECT 102.630 33.220 102.950 33.280 ;
        RECT 103.105 33.450 103.395 33.465 ;
        RECT 104.010 33.450 104.330 33.480 ;
        RECT 103.105 33.310 104.330 33.450 ;
        RECT 104.560 33.450 104.700 33.620 ;
        RECT 105.405 33.575 105.695 33.805 ;
        RECT 104.865 33.450 105.155 33.495 ;
        RECT 104.560 33.310 105.155 33.450 ;
        RECT 103.105 33.235 103.395 33.310 ;
        RECT 104.010 33.220 104.330 33.310 ;
        RECT 104.865 33.265 105.155 33.310 ;
        RECT 105.850 33.220 106.170 33.480 ;
        RECT 106.860 33.465 107.000 33.960 ;
        RECT 107.705 33.960 110.310 34.100 ;
        RECT 107.705 33.915 107.995 33.960 ;
        RECT 109.990 33.900 110.310 33.960 ;
        RECT 111.370 33.900 111.690 34.160 ;
        RECT 113.685 34.100 113.975 34.145 ;
        RECT 115.050 34.100 115.370 34.160 ;
        RECT 113.685 33.960 115.370 34.100 ;
        RECT 113.685 33.915 113.975 33.960 ;
        RECT 115.050 33.900 115.370 33.960 ;
        RECT 118.730 33.900 119.050 34.160 ;
        RECT 120.110 33.900 120.430 34.160 ;
        RECT 121.965 34.100 122.255 34.145 ;
        RECT 124.250 34.100 124.570 34.160 ;
        RECT 121.965 33.960 124.570 34.100 ;
        RECT 121.965 33.915 122.255 33.960 ;
        RECT 124.250 33.900 124.570 33.960 ;
        RECT 125.185 34.100 125.475 34.145 ;
        RECT 126.090 34.100 126.410 34.160 ;
        RECT 125.185 33.960 126.410 34.100 ;
        RECT 125.185 33.915 125.475 33.960 ;
        RECT 126.090 33.900 126.410 33.960 ;
        RECT 126.550 33.900 126.870 34.160 ;
        RECT 128.390 34.100 128.710 34.160 ;
        RECT 127.560 33.960 128.710 34.100 ;
        RECT 111.460 33.760 111.600 33.900 ;
        RECT 107.320 33.620 111.600 33.760 ;
        RECT 111.845 33.760 112.135 33.805 ;
        RECT 115.970 33.760 116.290 33.820 ;
        RECT 111.845 33.620 116.290 33.760 ;
        RECT 118.820 33.760 118.960 33.900 ;
        RECT 123.345 33.760 123.635 33.805 ;
        RECT 126.640 33.760 126.780 33.900 ;
        RECT 127.560 33.805 127.700 33.960 ;
        RECT 128.390 33.900 128.710 33.960 ;
        RECT 129.325 34.100 129.615 34.145 ;
        RECT 131.150 34.100 131.470 34.160 ;
        RECT 129.325 33.960 131.470 34.100 ;
        RECT 129.325 33.915 129.615 33.960 ;
        RECT 131.150 33.900 131.470 33.960 ;
        RECT 131.700 33.960 133.680 34.100 ;
        RECT 118.820 33.620 123.635 33.760 ;
        RECT 107.320 33.465 107.460 33.620 ;
        RECT 111.845 33.575 112.135 33.620 ;
        RECT 115.970 33.560 116.290 33.620 ;
        RECT 123.345 33.575 123.635 33.620 ;
        RECT 124.340 33.620 126.780 33.760 ;
        RECT 127.485 33.760 127.775 33.805 ;
        RECT 127.485 33.620 130.920 33.760 ;
        RECT 106.785 33.235 107.075 33.465 ;
        RECT 107.245 33.235 107.535 33.465 ;
        RECT 110.005 33.235 110.295 33.465 ;
        RECT 110.925 33.420 111.215 33.465 ;
        RECT 111.370 33.420 111.690 33.480 ;
        RECT 110.925 33.280 111.690 33.420 ;
        RECT 110.925 33.235 111.215 33.280 ;
        RECT 104.100 33.080 104.240 33.220 ;
        RECT 107.690 33.080 108.010 33.140 ;
        RECT 110.080 33.080 110.220 33.235 ;
        RECT 111.370 33.220 111.690 33.280 ;
        RECT 112.290 33.220 112.610 33.480 ;
        RECT 112.750 33.220 113.070 33.480 ;
        RECT 114.590 33.420 114.910 33.480 ;
        RECT 115.065 33.420 115.355 33.465 ;
        RECT 114.590 33.280 115.355 33.420 ;
        RECT 114.590 33.220 114.910 33.280 ;
        RECT 115.065 33.235 115.355 33.280 ;
        RECT 115.510 33.220 115.830 33.480 ;
        RECT 117.810 33.220 118.130 33.480 ;
        RECT 119.205 33.420 119.495 33.465 ;
        RECT 118.360 33.280 119.495 33.420 ;
        RECT 114.145 33.080 114.435 33.125 ;
        RECT 104.100 32.940 110.220 33.080 ;
        RECT 110.540 32.940 114.435 33.080 ;
        RECT 115.600 33.080 115.740 33.220 ;
        RECT 118.360 33.080 118.500 33.280 ;
        RECT 119.205 33.235 119.495 33.280 ;
        RECT 122.425 33.235 122.715 33.465 ;
        RECT 115.600 32.940 118.500 33.080 ;
        RECT 118.745 33.080 119.035 33.125 ;
        RECT 122.500 33.080 122.640 33.235 ;
        RECT 122.870 33.220 123.190 33.480 ;
        RECT 124.340 33.465 124.480 33.620 ;
        RECT 127.485 33.575 127.775 33.620 ;
        RECT 124.265 33.235 124.555 33.465 ;
        RECT 126.565 33.420 126.855 33.465 ;
        RECT 127.010 33.420 127.330 33.480 ;
        RECT 126.565 33.280 127.330 33.420 ;
        RECT 126.565 33.235 126.855 33.280 ;
        RECT 127.010 33.220 127.330 33.280 ;
        RECT 127.930 33.220 128.250 33.480 ;
        RECT 128.405 33.420 128.695 33.465 ;
        RECT 130.230 33.420 130.550 33.480 ;
        RECT 128.405 33.280 130.550 33.420 ;
        RECT 128.405 33.235 128.695 33.280 ;
        RECT 128.480 33.080 128.620 33.235 ;
        RECT 130.230 33.220 130.550 33.280 ;
        RECT 118.745 32.940 128.620 33.080 ;
        RECT 130.780 33.080 130.920 33.620 ;
        RECT 131.165 33.420 131.455 33.465 ;
        RECT 131.700 33.420 131.840 33.960 ;
        RECT 132.070 33.560 132.390 33.820 ;
        RECT 133.540 33.760 133.680 33.960 ;
        RECT 133.910 33.900 134.230 34.160 ;
        RECT 146.330 34.100 146.650 34.160 ;
        RECT 146.805 34.100 147.095 34.145 ;
        RECT 146.330 33.960 147.095 34.100 ;
        RECT 146.330 33.900 146.650 33.960 ;
        RECT 146.805 33.915 147.095 33.960 ;
        RECT 148.185 34.100 148.475 34.145 ;
        RECT 149.090 34.100 149.410 34.160 ;
        RECT 148.185 33.960 149.410 34.100 ;
        RECT 148.185 33.915 148.475 33.960 ;
        RECT 149.090 33.900 149.410 33.960 ;
        RECT 149.550 33.900 149.870 34.160 ;
        RECT 137.590 33.760 137.910 33.820 ;
        RECT 133.540 33.620 134.600 33.760 ;
        RECT 131.165 33.280 131.840 33.420 ;
        RECT 132.160 33.420 132.300 33.560 ;
        RECT 134.460 33.480 134.600 33.620 ;
        RECT 137.590 33.620 147.480 33.760 ;
        RECT 137.590 33.560 137.910 33.620 ;
        RECT 132.545 33.420 132.835 33.465 ;
        RECT 132.160 33.280 132.835 33.420 ;
        RECT 131.165 33.235 131.455 33.280 ;
        RECT 132.545 33.235 132.835 33.280 ;
        RECT 133.005 33.420 133.295 33.465 ;
        RECT 133.005 33.280 133.405 33.420 ;
        RECT 133.005 33.235 133.295 33.280 ;
        RECT 133.080 33.080 133.220 33.235 ;
        RECT 134.370 33.220 134.690 33.480 ;
        RECT 145.870 33.420 146.190 33.480 ;
        RECT 147.340 33.465 147.480 33.620 ;
        RECT 146.345 33.420 146.635 33.465 ;
        RECT 145.870 33.280 146.635 33.420 ;
        RECT 145.870 33.220 146.190 33.280 ;
        RECT 146.345 33.235 146.635 33.280 ;
        RECT 147.265 33.235 147.555 33.465 ;
        RECT 147.725 33.420 148.015 33.465 ;
        RECT 149.640 33.420 149.780 33.900 ;
        RECT 147.725 33.280 149.780 33.420 ;
        RECT 150.485 33.420 150.775 33.465 ;
        RECT 152.770 33.420 153.090 33.480 ;
        RECT 150.485 33.280 153.090 33.420 ;
        RECT 147.725 33.235 148.015 33.280 ;
        RECT 150.485 33.235 150.775 33.280 ;
        RECT 152.770 33.220 153.090 33.280 ;
        RECT 137.590 33.080 137.910 33.140 ;
        RECT 130.780 32.940 137.910 33.080 ;
        RECT 107.690 32.880 108.010 32.940 ;
        RECT 105.390 32.740 105.710 32.800 ;
        RECT 102.720 32.600 105.710 32.740 ;
        RECT 99.425 32.400 99.715 32.445 ;
        RECT 102.170 32.400 102.490 32.460 ;
        RECT 102.720 32.445 102.860 32.600 ;
        RECT 105.390 32.540 105.710 32.600 ;
        RECT 105.850 32.740 106.170 32.800 ;
        RECT 108.165 32.740 108.455 32.785 ;
        RECT 105.850 32.600 108.455 32.740 ;
        RECT 105.850 32.540 106.170 32.600 ;
        RECT 108.165 32.555 108.455 32.600 ;
        RECT 109.530 32.740 109.850 32.800 ;
        RECT 110.540 32.740 110.680 32.940 ;
        RECT 114.145 32.895 114.435 32.940 ;
        RECT 118.745 32.895 119.035 32.940 ;
        RECT 137.590 32.880 137.910 32.940 ;
        RECT 139.890 33.080 140.210 33.140 ;
        RECT 139.890 32.940 149.780 33.080 ;
        RECT 139.890 32.880 140.210 32.940 ;
        RECT 109.530 32.600 110.680 32.740 ;
        RECT 127.470 32.740 127.790 32.800 ;
        RECT 131.625 32.740 131.915 32.785 ;
        RECT 140.810 32.740 141.130 32.800 ;
        RECT 149.640 32.785 149.780 32.940 ;
        RECT 127.470 32.600 141.130 32.740 ;
        RECT 109.530 32.540 109.850 32.600 ;
        RECT 127.470 32.540 127.790 32.600 ;
        RECT 131.625 32.555 131.915 32.600 ;
        RECT 140.810 32.540 141.130 32.600 ;
        RECT 149.565 32.555 149.855 32.785 ;
        RECT 99.425 32.260 102.490 32.400 ;
        RECT 99.425 32.215 99.715 32.260 ;
        RECT 102.170 32.200 102.490 32.260 ;
        RECT 102.645 32.215 102.935 32.445 ;
        RECT 104.025 32.400 104.315 32.445 ;
        RECT 110.910 32.400 111.230 32.460 ;
        RECT 104.025 32.260 111.230 32.400 ;
        RECT 104.025 32.215 104.315 32.260 ;
        RECT 110.910 32.200 111.230 32.260 ;
        RECT 111.370 32.400 111.690 32.460 ;
        RECT 117.825 32.400 118.115 32.445 ;
        RECT 111.370 32.260 118.115 32.400 ;
        RECT 111.370 32.200 111.690 32.260 ;
        RECT 117.825 32.215 118.115 32.260 ;
        RECT 153.860 32.060 154.340 34.170 ;
        RECT 91.060 31.580 154.340 32.060 ;
        RECT 93.430 31.180 93.750 31.440 ;
        RECT 99.425 31.380 99.715 31.425 ;
        RECT 99.870 31.380 100.190 31.440 ;
        RECT 99.425 31.240 100.190 31.380 ;
        RECT 99.425 31.195 99.715 31.240 ;
        RECT 99.870 31.180 100.190 31.240 ;
        RECT 107.245 31.380 107.535 31.425 ;
        RECT 107.690 31.380 108.010 31.440 ;
        RECT 111.370 31.380 111.690 31.440 ;
        RECT 107.245 31.240 111.690 31.380 ;
        RECT 107.245 31.195 107.535 31.240 ;
        RECT 107.690 31.180 108.010 31.240 ;
        RECT 111.370 31.180 111.690 31.240 ;
        RECT 115.065 31.380 115.355 31.425 ;
        RECT 115.510 31.380 115.830 31.440 ;
        RECT 115.065 31.240 115.830 31.380 ;
        RECT 115.065 31.195 115.355 31.240 ;
        RECT 115.510 31.180 115.830 31.240 ;
        RECT 117.810 31.180 118.130 31.440 ;
        RECT 130.230 31.180 130.550 31.440 ;
        RECT 137.590 31.180 137.910 31.440 ;
        RECT 149.565 31.380 149.855 31.425 ;
        RECT 150.930 31.380 151.250 31.440 ;
        RECT 149.565 31.240 151.250 31.380 ;
        RECT 149.565 31.195 149.855 31.240 ;
        RECT 150.930 31.180 151.250 31.240 ;
        RECT 117.900 31.040 118.040 31.180 ;
        RECT 121.965 31.040 122.255 31.085 ;
        RECT 117.900 30.900 122.255 31.040 ;
        RECT 90.210 30.360 90.530 30.420 ;
        RECT 92.525 30.360 92.815 30.405 ;
        RECT 90.210 30.220 92.815 30.360 ;
        RECT 90.210 30.160 90.530 30.220 ;
        RECT 92.525 30.175 92.815 30.220 ;
        RECT 98.490 30.160 98.810 30.420 ;
        RECT 106.310 30.160 106.630 30.420 ;
        RECT 114.130 30.160 114.450 30.420 ;
        RECT 115.970 30.360 116.290 30.420 ;
        RECT 119.740 30.405 119.880 30.900 ;
        RECT 121.965 30.855 122.255 30.900 ;
        RECT 140.810 30.700 141.130 30.760 ;
        RECT 144.505 30.700 144.795 30.745 ;
        RECT 140.810 30.560 144.795 30.700 ;
        RECT 140.810 30.500 141.130 30.560 ;
        RECT 144.505 30.515 144.795 30.560 ;
        RECT 119.205 30.360 119.495 30.405 ;
        RECT 115.970 30.220 119.495 30.360 ;
        RECT 115.970 30.160 116.290 30.220 ;
        RECT 119.205 30.175 119.495 30.220 ;
        RECT 119.665 30.175 119.955 30.405 ;
        RECT 121.490 30.360 121.810 30.420 ;
        RECT 122.885 30.360 123.175 30.405 ;
        RECT 121.490 30.220 123.175 30.360 ;
        RECT 121.490 30.160 121.810 30.220 ;
        RECT 122.885 30.175 123.175 30.220 ;
        RECT 129.310 30.360 129.630 30.420 ;
        RECT 131.165 30.360 131.455 30.405 ;
        RECT 129.310 30.220 131.455 30.360 ;
        RECT 129.310 30.160 129.630 30.220 ;
        RECT 131.165 30.175 131.455 30.220 ;
        RECT 137.130 30.360 137.450 30.420 ;
        RECT 138.525 30.360 138.815 30.405 ;
        RECT 137.130 30.220 138.815 30.360 ;
        RECT 137.130 30.160 137.450 30.220 ;
        RECT 138.525 30.175 138.815 30.220 ;
        RECT 143.125 30.175 143.415 30.405 ;
        RECT 143.200 30.020 143.340 30.175 ;
        RECT 144.950 30.020 145.270 30.080 ;
        RECT 143.200 29.880 145.270 30.020 ;
        RECT 144.950 29.820 145.270 29.880 ;
        RECT 150.025 30.020 150.315 30.065 ;
        RECT 151.850 30.020 152.170 30.080 ;
        RECT 150.025 29.880 152.170 30.020 ;
        RECT 150.025 29.835 150.315 29.880 ;
        RECT 151.850 29.820 152.170 29.880 ;
        RECT 88.980 28.860 152.240 29.340 ;
        RECT 1.000 24.610 2.510 25.490 ;
        RECT 1.000 24.130 57.585 24.610 ;
        RECT 59.105 24.375 59.355 26.480 ;
        RECT 61.215 24.610 61.695 24.615 ;
        RECT 153.860 24.610 154.340 31.580 ;
        RECT 61.215 24.130 154.340 24.610 ;
        RECT 1.000 23.170 2.510 24.130 ;
        RECT 57.095 23.190 57.575 24.130 ;
        RECT 61.215 23.190 61.695 24.130 ;
        RECT 57.095 22.710 61.695 23.190 ;
        RECT 6.070 19.805 6.320 21.910 ;
        RECT 59.010 20.540 59.440 20.940 ;
        RECT 6.070 16.650 6.320 18.755 ;
        RECT 8.230 15.990 10.045 18.735 ;
        RECT 59.110 10.455 59.360 12.560 ;
        RECT 53.125 7.780 54.035 8.675 ;
        RECT 59.110 7.800 59.360 9.905 ;
        RECT 82.960 7.520 83.920 8.410 ;
      LAYER via ;
        RECT 84.955 222.590 85.215 222.850 ;
        RECT 84.950 200.305 85.210 200.565 ;
        RECT 1.495 194.185 1.995 194.685 ;
        RECT 76.515 194.300 76.775 194.560 ;
        RECT 76.835 194.300 77.095 194.560 ;
        RECT 77.155 194.300 77.415 194.560 ;
        RECT 77.475 194.300 77.735 194.560 ;
        RECT 77.795 194.300 78.055 194.560 ;
        RECT 88.590 194.300 88.850 194.560 ;
        RECT 88.910 194.300 89.170 194.560 ;
        RECT 89.230 194.300 89.490 194.560 ;
        RECT 89.550 194.300 89.810 194.560 ;
        RECT 89.870 194.300 90.130 194.560 ;
        RECT 100.665 194.300 100.925 194.560 ;
        RECT 100.985 194.300 101.245 194.560 ;
        RECT 101.305 194.300 101.565 194.560 ;
        RECT 101.625 194.300 101.885 194.560 ;
        RECT 101.945 194.300 102.205 194.560 ;
        RECT 112.740 194.300 113.000 194.560 ;
        RECT 113.060 194.300 113.320 194.560 ;
        RECT 113.380 194.300 113.640 194.560 ;
        RECT 113.700 194.300 113.960 194.560 ;
        RECT 114.020 194.300 114.280 194.560 ;
        RECT 80.550 193.790 80.810 194.050 ;
        RECT 110.450 193.790 110.710 194.050 ;
        RECT 86.990 192.770 87.250 193.030 ;
        RECT 81.470 192.430 81.730 192.690 ;
        RECT 100.330 192.430 100.590 192.690 ;
        RECT 102.630 192.430 102.890 192.690 ;
        RECT 111.370 192.430 111.630 192.690 ;
        RECT 82.390 192.090 82.650 192.350 ;
        RECT 106.770 192.090 107.030 192.350 ;
        RECT 79.815 191.580 80.075 191.840 ;
        RECT 80.135 191.580 80.395 191.840 ;
        RECT 80.455 191.580 80.715 191.840 ;
        RECT 80.775 191.580 81.035 191.840 ;
        RECT 81.095 191.580 81.355 191.840 ;
        RECT 91.890 191.580 92.150 191.840 ;
        RECT 92.210 191.580 92.470 191.840 ;
        RECT 92.530 191.580 92.790 191.840 ;
        RECT 92.850 191.580 93.110 191.840 ;
        RECT 93.170 191.580 93.430 191.840 ;
        RECT 103.965 191.580 104.225 191.840 ;
        RECT 104.285 191.580 104.545 191.840 ;
        RECT 104.605 191.580 104.865 191.840 ;
        RECT 104.925 191.580 105.185 191.840 ;
        RECT 105.245 191.580 105.505 191.840 ;
        RECT 116.040 191.580 116.300 191.840 ;
        RECT 116.360 191.580 116.620 191.840 ;
        RECT 116.680 191.580 116.940 191.840 ;
        RECT 117.000 191.580 117.260 191.840 ;
        RECT 117.320 191.580 117.580 191.840 ;
        RECT 81.470 191.070 81.730 191.330 ;
        RECT 70.430 190.390 70.690 190.650 ;
        RECT 81.010 190.390 81.270 190.650 ;
        RECT 82.850 190.390 83.110 190.650 ;
        RECT 106.310 191.070 106.570 191.330 ;
        RECT 111.370 191.070 111.630 191.330 ;
        RECT 107.690 190.730 107.950 190.990 ;
        RECT 87.910 190.050 88.170 190.310 ;
        RECT 100.330 190.390 100.590 190.650 ;
        RECT 103.090 190.390 103.350 190.650 ;
        RECT 104.470 190.390 104.730 190.650 ;
        RECT 83.770 189.710 84.030 189.970 ;
        RECT 73.650 189.370 73.910 189.630 ;
        RECT 84.230 189.370 84.490 189.630 ;
        RECT 86.990 189.370 87.250 189.630 ;
        RECT 94.810 190.050 95.070 190.310 ;
        RECT 104.010 190.050 104.270 190.310 ;
        RECT 93.890 189.370 94.150 189.630 ;
        RECT 94.350 189.370 94.610 189.630 ;
        RECT 103.550 189.370 103.810 189.630 ;
        RECT 109.070 190.390 109.330 190.650 ;
        RECT 120.110 189.710 120.370 189.970 ;
        RECT 111.830 189.370 112.090 189.630 ;
        RECT 76.515 188.860 76.775 189.120 ;
        RECT 76.835 188.860 77.095 189.120 ;
        RECT 77.155 188.860 77.415 189.120 ;
        RECT 77.475 188.860 77.735 189.120 ;
        RECT 77.795 188.860 78.055 189.120 ;
        RECT 88.590 188.860 88.850 189.120 ;
        RECT 88.910 188.860 89.170 189.120 ;
        RECT 89.230 188.860 89.490 189.120 ;
        RECT 89.550 188.860 89.810 189.120 ;
        RECT 89.870 188.860 90.130 189.120 ;
        RECT 100.665 188.860 100.925 189.120 ;
        RECT 100.985 188.860 101.245 189.120 ;
        RECT 101.305 188.860 101.565 189.120 ;
        RECT 101.625 188.860 101.885 189.120 ;
        RECT 101.945 188.860 102.205 189.120 ;
        RECT 112.740 188.860 113.000 189.120 ;
        RECT 113.060 188.860 113.320 189.120 ;
        RECT 113.380 188.860 113.640 189.120 ;
        RECT 113.700 188.860 113.960 189.120 ;
        RECT 114.020 188.860 114.280 189.120 ;
        RECT 73.650 188.350 73.910 188.610 ;
        RECT 82.390 188.350 82.650 188.610 ;
        RECT 82.850 188.350 83.110 188.610 ;
        RECT 94.350 188.350 94.610 188.610 ;
        RECT 104.010 188.350 104.270 188.610 ;
        RECT 107.690 188.350 107.950 188.610 ;
        RECT 106.310 188.010 106.570 188.270 ;
        RECT 83.770 187.330 84.030 187.590 ;
        RECT 93.890 187.670 94.150 187.930 ;
        RECT 104.470 187.670 104.730 187.930 ;
        RECT 94.810 187.330 95.070 187.590 ;
        RECT 84.230 186.990 84.490 187.250 ;
        RECT 89.290 186.990 89.550 187.250 ;
        RECT 85.150 186.650 85.410 186.910 ;
        RECT 99.870 187.330 100.130 187.590 ;
        RECT 98.490 186.990 98.750 187.250 ;
        RECT 101.250 186.990 101.510 187.250 ;
        RECT 106.770 187.330 107.030 187.590 ;
        RECT 108.150 187.670 108.410 187.930 ;
        RECT 111.830 187.670 112.090 187.930 ;
        RECT 119.190 188.350 119.450 188.610 ;
        RECT 102.630 186.650 102.890 186.910 ;
        RECT 113.210 186.650 113.470 186.910 ;
        RECT 79.815 186.140 80.075 186.400 ;
        RECT 80.135 186.140 80.395 186.400 ;
        RECT 80.455 186.140 80.715 186.400 ;
        RECT 80.775 186.140 81.035 186.400 ;
        RECT 81.095 186.140 81.355 186.400 ;
        RECT 91.890 186.140 92.150 186.400 ;
        RECT 92.210 186.140 92.470 186.400 ;
        RECT 92.530 186.140 92.790 186.400 ;
        RECT 92.850 186.140 93.110 186.400 ;
        RECT 93.170 186.140 93.430 186.400 ;
        RECT 103.965 186.140 104.225 186.400 ;
        RECT 104.285 186.140 104.545 186.400 ;
        RECT 104.605 186.140 104.865 186.400 ;
        RECT 104.925 186.140 105.185 186.400 ;
        RECT 105.245 186.140 105.505 186.400 ;
        RECT 116.040 186.140 116.300 186.400 ;
        RECT 116.360 186.140 116.620 186.400 ;
        RECT 116.680 186.140 116.940 186.400 ;
        RECT 117.000 186.140 117.260 186.400 ;
        RECT 117.320 186.140 117.580 186.400 ;
        RECT 79.170 185.630 79.430 185.890 ;
        RECT 83.770 185.630 84.030 185.890 ;
        RECT 89.290 185.630 89.550 185.890 ;
        RECT 98.490 185.630 98.750 185.890 ;
        RECT 98.950 185.630 99.210 185.890 ;
        RECT 103.550 185.630 103.810 185.890 ;
        RECT 106.310 185.630 106.570 185.890 ;
        RECT 108.150 185.630 108.410 185.890 ;
        RECT 85.150 184.950 85.410 185.210 ;
        RECT 94.350 184.950 94.610 185.210 ;
        RECT 101.250 184.950 101.510 185.210 ;
        RECT 102.630 184.950 102.890 185.210 ;
        RECT 103.090 184.950 103.350 185.210 ;
        RECT 113.210 185.290 113.470 185.550 ;
        RECT 87.910 184.610 88.170 184.870 ;
        RECT 91.130 184.610 91.390 184.870 ;
        RECT 100.330 184.610 100.590 184.870 ;
        RECT 106.310 184.610 106.570 184.870 ;
        RECT 83.770 183.930 84.030 184.190 ;
        RECT 86.990 184.270 87.250 184.530 ;
        RECT 92.970 184.270 93.230 184.530 ;
        RECT 110.910 184.610 111.170 184.870 ;
        RECT 95.730 183.930 95.990 184.190 ;
        RECT 106.770 183.930 107.030 184.190 ;
        RECT 76.515 183.420 76.775 183.680 ;
        RECT 76.835 183.420 77.095 183.680 ;
        RECT 77.155 183.420 77.415 183.680 ;
        RECT 77.475 183.420 77.735 183.680 ;
        RECT 77.795 183.420 78.055 183.680 ;
        RECT 88.590 183.420 88.850 183.680 ;
        RECT 88.910 183.420 89.170 183.680 ;
        RECT 89.230 183.420 89.490 183.680 ;
        RECT 89.550 183.420 89.810 183.680 ;
        RECT 89.870 183.420 90.130 183.680 ;
        RECT 100.665 183.420 100.925 183.680 ;
        RECT 100.985 183.420 101.245 183.680 ;
        RECT 101.305 183.420 101.565 183.680 ;
        RECT 101.625 183.420 101.885 183.680 ;
        RECT 101.945 183.420 102.205 183.680 ;
        RECT 112.740 183.420 113.000 183.680 ;
        RECT 113.060 183.420 113.320 183.680 ;
        RECT 113.380 183.420 113.640 183.680 ;
        RECT 113.700 183.420 113.960 183.680 ;
        RECT 114.020 183.420 114.280 183.680 ;
        RECT 83.770 182.910 84.030 183.170 ;
        RECT 87.910 182.910 88.170 183.170 ;
        RECT 91.130 182.910 91.390 183.170 ;
        RECT 94.350 182.910 94.610 183.170 ;
        RECT 92.970 181.890 93.230 182.150 ;
        RECT 95.730 181.890 95.990 182.150 ;
        RECT 98.950 182.570 99.210 182.830 ;
        RECT 93.890 181.550 94.150 181.810 ;
        RECT 102.630 181.550 102.890 181.810 ;
        RECT 100.330 181.210 100.590 181.470 ;
        RECT 105.850 181.550 106.110 181.810 ;
        RECT 115.050 181.550 115.310 181.810 ;
        RECT 106.310 181.210 106.570 181.470 ;
        RECT 111.830 181.210 112.090 181.470 ;
        RECT 79.815 180.700 80.075 180.960 ;
        RECT 80.135 180.700 80.395 180.960 ;
        RECT 80.455 180.700 80.715 180.960 ;
        RECT 80.775 180.700 81.035 180.960 ;
        RECT 81.095 180.700 81.355 180.960 ;
        RECT 91.890 180.700 92.150 180.960 ;
        RECT 92.210 180.700 92.470 180.960 ;
        RECT 92.530 180.700 92.790 180.960 ;
        RECT 92.850 180.700 93.110 180.960 ;
        RECT 93.170 180.700 93.430 180.960 ;
        RECT 103.965 180.700 104.225 180.960 ;
        RECT 104.285 180.700 104.545 180.960 ;
        RECT 104.605 180.700 104.865 180.960 ;
        RECT 104.925 180.700 105.185 180.960 ;
        RECT 105.245 180.700 105.505 180.960 ;
        RECT 116.040 180.700 116.300 180.960 ;
        RECT 116.360 180.700 116.620 180.960 ;
        RECT 116.680 180.700 116.940 180.960 ;
        RECT 117.000 180.700 117.260 180.960 ;
        RECT 117.320 180.700 117.580 180.960 ;
        RECT 99.410 180.190 99.670 180.450 ;
        RECT 107.690 180.190 107.950 180.450 ;
        RECT 110.910 180.190 111.170 180.450 ;
        RECT 73.650 179.510 73.910 179.770 ;
        RECT 82.390 179.510 82.650 179.770 ;
        RECT 75.030 179.170 75.290 179.430 ;
        RECT 99.870 179.850 100.130 180.110 ;
        RECT 100.330 179.510 100.590 179.770 ;
        RECT 105.850 179.510 106.110 179.770 ;
        RECT 106.770 179.510 107.030 179.770 ;
        RECT 85.610 178.830 85.870 179.090 ;
        RECT 85.150 178.490 85.410 178.750 ;
        RECT 97.110 178.490 97.370 178.750 ;
        RECT 112.290 178.490 112.550 178.750 ;
        RECT 76.515 177.980 76.775 178.240 ;
        RECT 76.835 177.980 77.095 178.240 ;
        RECT 77.155 177.980 77.415 178.240 ;
        RECT 77.475 177.980 77.735 178.240 ;
        RECT 77.795 177.980 78.055 178.240 ;
        RECT 88.590 177.980 88.850 178.240 ;
        RECT 88.910 177.980 89.170 178.240 ;
        RECT 89.230 177.980 89.490 178.240 ;
        RECT 89.550 177.980 89.810 178.240 ;
        RECT 89.870 177.980 90.130 178.240 ;
        RECT 100.665 177.980 100.925 178.240 ;
        RECT 100.985 177.980 101.245 178.240 ;
        RECT 101.305 177.980 101.565 178.240 ;
        RECT 101.625 177.980 101.885 178.240 ;
        RECT 101.945 177.980 102.205 178.240 ;
        RECT 112.740 177.980 113.000 178.240 ;
        RECT 113.060 177.980 113.320 178.240 ;
        RECT 113.380 177.980 113.640 178.240 ;
        RECT 113.700 177.980 113.960 178.240 ;
        RECT 114.020 177.980 114.280 178.240 ;
        RECT 75.030 177.470 75.290 177.730 ;
        RECT 99.870 177.470 100.130 177.730 ;
        RECT 96.190 177.130 96.450 177.390 ;
        RECT 103.090 177.470 103.350 177.730 ;
        RECT 115.050 177.470 115.310 177.730 ;
        RECT 81.470 176.790 81.730 177.050 ;
        RECT 85.150 176.790 85.410 177.050 ;
        RECT 111.370 176.790 111.630 177.050 ;
        RECT 82.850 176.450 83.110 176.710 ;
        RECT 97.110 176.450 97.370 176.710 ;
        RECT 103.550 176.450 103.810 176.710 ;
        RECT 108.610 176.450 108.870 176.710 ;
        RECT 112.290 176.450 112.550 176.710 ;
        RECT 118.730 176.790 118.990 177.050 ;
        RECT 83.770 176.110 84.030 176.370 ;
        RECT 96.650 176.110 96.910 176.370 ;
        RECT 105.850 175.770 106.110 176.030 ;
        RECT 107.230 175.770 107.490 176.030 ;
        RECT 114.590 175.770 114.850 176.030 ;
        RECT 115.050 175.770 115.310 176.030 ;
        RECT 115.510 175.770 115.770 176.030 ;
        RECT 117.810 175.770 118.070 176.030 ;
        RECT 79.815 175.260 80.075 175.520 ;
        RECT 80.135 175.260 80.395 175.520 ;
        RECT 80.455 175.260 80.715 175.520 ;
        RECT 80.775 175.260 81.035 175.520 ;
        RECT 81.095 175.260 81.355 175.520 ;
        RECT 91.890 175.260 92.150 175.520 ;
        RECT 92.210 175.260 92.470 175.520 ;
        RECT 92.530 175.260 92.790 175.520 ;
        RECT 92.850 175.260 93.110 175.520 ;
        RECT 93.170 175.260 93.430 175.520 ;
        RECT 103.965 175.260 104.225 175.520 ;
        RECT 104.285 175.260 104.545 175.520 ;
        RECT 104.605 175.260 104.865 175.520 ;
        RECT 104.925 175.260 105.185 175.520 ;
        RECT 105.245 175.260 105.505 175.520 ;
        RECT 116.040 175.260 116.300 175.520 ;
        RECT 116.360 175.260 116.620 175.520 ;
        RECT 116.680 175.260 116.940 175.520 ;
        RECT 117.000 175.260 117.260 175.520 ;
        RECT 117.320 175.260 117.580 175.520 ;
        RECT 73.650 174.070 73.910 174.330 ;
        RECT 79.170 174.750 79.430 175.010 ;
        RECT 75.490 173.730 75.750 173.990 ;
        RECT 82.390 174.070 82.650 174.330 ;
        RECT 99.870 174.750 100.130 175.010 ;
        RECT 103.550 174.750 103.810 175.010 ;
        RECT 107.230 174.750 107.490 175.010 ;
        RECT 108.610 174.750 108.870 175.010 ;
        RECT 111.830 174.750 112.090 175.010 ;
        RECT 81.470 173.730 81.730 173.990 ;
        RECT 82.850 173.050 83.110 173.310 ;
        RECT 93.890 174.070 94.150 174.330 ;
        RECT 97.110 174.070 97.370 174.330 ;
        RECT 106.310 174.410 106.570 174.670 ;
        RECT 96.190 173.730 96.450 173.990 ;
        RECT 107.690 174.070 107.950 174.330 ;
        RECT 117.350 174.070 117.610 174.330 ;
        RECT 117.810 174.070 118.070 174.330 ;
        RECT 108.610 173.730 108.870 173.990 ;
        RECT 111.370 173.730 111.630 173.990 ;
        RECT 115.050 173.730 115.310 173.990 ;
        RECT 93.430 173.050 93.690 173.310 ;
        RECT 115.050 173.050 115.310 173.310 ;
        RECT 118.270 173.050 118.530 173.310 ;
        RECT 76.515 172.540 76.775 172.800 ;
        RECT 76.835 172.540 77.095 172.800 ;
        RECT 77.155 172.540 77.415 172.800 ;
        RECT 77.475 172.540 77.735 172.800 ;
        RECT 77.795 172.540 78.055 172.800 ;
        RECT 88.590 172.540 88.850 172.800 ;
        RECT 88.910 172.540 89.170 172.800 ;
        RECT 89.230 172.540 89.490 172.800 ;
        RECT 89.550 172.540 89.810 172.800 ;
        RECT 89.870 172.540 90.130 172.800 ;
        RECT 100.665 172.540 100.925 172.800 ;
        RECT 100.985 172.540 101.245 172.800 ;
        RECT 101.305 172.540 101.565 172.800 ;
        RECT 101.625 172.540 101.885 172.800 ;
        RECT 101.945 172.540 102.205 172.800 ;
        RECT 112.740 172.540 113.000 172.800 ;
        RECT 113.060 172.540 113.320 172.800 ;
        RECT 113.380 172.540 113.640 172.800 ;
        RECT 113.700 172.540 113.960 172.800 ;
        RECT 114.020 172.540 114.280 172.800 ;
        RECT 75.490 172.030 75.750 172.290 ;
        RECT 83.770 172.030 84.030 172.290 ;
        RECT 108.610 172.030 108.870 172.290 ;
        RECT 75.030 171.350 75.290 171.610 ;
        RECT 81.470 171.350 81.730 171.610 ;
        RECT 82.390 171.350 82.650 171.610 ;
        RECT 93.430 171.350 93.690 171.610 ;
        RECT 117.350 171.690 117.610 171.950 ;
        RECT 115.050 171.350 115.310 171.610 ;
        RECT 82.850 171.010 83.110 171.270 ;
        RECT 86.530 170.670 86.790 170.930 ;
        RECT 103.090 170.670 103.350 170.930 ;
        RECT 81.470 170.330 81.730 170.590 ;
        RECT 96.650 170.330 96.910 170.590 ;
        RECT 108.150 170.330 108.410 170.590 ;
        RECT 114.130 170.330 114.390 170.590 ;
        RECT 79.815 169.820 80.075 170.080 ;
        RECT 80.135 169.820 80.395 170.080 ;
        RECT 80.455 169.820 80.715 170.080 ;
        RECT 80.775 169.820 81.035 170.080 ;
        RECT 81.095 169.820 81.355 170.080 ;
        RECT 91.890 169.820 92.150 170.080 ;
        RECT 92.210 169.820 92.470 170.080 ;
        RECT 92.530 169.820 92.790 170.080 ;
        RECT 92.850 169.820 93.110 170.080 ;
        RECT 93.170 169.820 93.430 170.080 ;
        RECT 103.965 169.820 104.225 170.080 ;
        RECT 104.285 169.820 104.545 170.080 ;
        RECT 104.605 169.820 104.865 170.080 ;
        RECT 104.925 169.820 105.185 170.080 ;
        RECT 105.245 169.820 105.505 170.080 ;
        RECT 116.040 169.820 116.300 170.080 ;
        RECT 116.360 169.820 116.620 170.080 ;
        RECT 116.680 169.820 116.940 170.080 ;
        RECT 117.000 169.820 117.260 170.080 ;
        RECT 117.320 169.820 117.580 170.080 ;
        RECT 103.090 169.310 103.350 169.570 ;
        RECT 105.850 169.310 106.110 169.570 ;
        RECT 85.610 168.630 85.870 168.890 ;
        RECT 90.210 168.630 90.470 168.890 ;
        RECT 93.890 168.630 94.150 168.890 ;
        RECT 114.130 169.310 114.390 169.570 ;
        RECT 117.810 169.310 118.070 169.570 ;
        RECT 107.690 168.630 107.950 168.890 ;
        RECT 82.390 168.290 82.650 168.550 ;
        RECT 83.770 168.290 84.030 168.550 ;
        RECT 93.890 167.610 94.150 167.870 ;
        RECT 94.810 167.610 95.070 167.870 ;
        RECT 95.730 167.610 95.990 167.870 ;
        RECT 108.150 167.610 108.410 167.870 ;
        RECT 76.515 167.100 76.775 167.360 ;
        RECT 76.835 167.100 77.095 167.360 ;
        RECT 77.155 167.100 77.415 167.360 ;
        RECT 77.475 167.100 77.735 167.360 ;
        RECT 77.795 167.100 78.055 167.360 ;
        RECT 88.590 167.100 88.850 167.360 ;
        RECT 88.910 167.100 89.170 167.360 ;
        RECT 89.230 167.100 89.490 167.360 ;
        RECT 89.550 167.100 89.810 167.360 ;
        RECT 89.870 167.100 90.130 167.360 ;
        RECT 100.665 167.100 100.925 167.360 ;
        RECT 100.985 167.100 101.245 167.360 ;
        RECT 101.305 167.100 101.565 167.360 ;
        RECT 101.625 167.100 101.885 167.360 ;
        RECT 101.945 167.100 102.205 167.360 ;
        RECT 112.740 167.100 113.000 167.360 ;
        RECT 113.060 167.100 113.320 167.360 ;
        RECT 113.380 167.100 113.640 167.360 ;
        RECT 113.700 167.100 113.960 167.360 ;
        RECT 114.020 167.100 114.280 167.360 ;
        RECT 75.030 166.590 75.290 166.850 ;
        RECT 106.310 166.590 106.570 166.850 ;
        RECT 115.510 166.590 115.770 166.850 ;
        RECT 81.470 165.910 81.730 166.170 ;
        RECT 82.390 165.910 82.650 166.170 ;
        RECT 94.810 165.910 95.070 166.170 ;
        RECT 81.010 165.570 81.270 165.830 ;
        RECT 85.610 165.570 85.870 165.830 ;
        RECT 114.590 165.570 114.850 165.830 ;
        RECT 118.270 165.230 118.530 165.490 ;
        RECT 76.870 164.890 77.130 165.150 ;
        RECT 89.290 164.890 89.550 165.150 ;
        RECT 90.210 164.890 90.470 165.150 ;
        RECT 93.890 164.890 94.150 165.150 ;
        RECT 95.730 164.890 95.990 165.150 ;
        RECT 106.770 164.890 107.030 165.150 ;
        RECT 110.450 164.890 110.710 165.150 ;
        RECT 111.830 164.890 112.090 165.150 ;
        RECT 115.050 164.890 115.310 165.150 ;
        RECT 79.815 164.380 80.075 164.640 ;
        RECT 80.135 164.380 80.395 164.640 ;
        RECT 80.455 164.380 80.715 164.640 ;
        RECT 80.775 164.380 81.035 164.640 ;
        RECT 81.095 164.380 81.355 164.640 ;
        RECT 91.890 164.380 92.150 164.640 ;
        RECT 92.210 164.380 92.470 164.640 ;
        RECT 92.530 164.380 92.790 164.640 ;
        RECT 92.850 164.380 93.110 164.640 ;
        RECT 93.170 164.380 93.430 164.640 ;
        RECT 103.965 164.380 104.225 164.640 ;
        RECT 104.285 164.380 104.545 164.640 ;
        RECT 104.605 164.380 104.865 164.640 ;
        RECT 104.925 164.380 105.185 164.640 ;
        RECT 105.245 164.380 105.505 164.640 ;
        RECT 116.040 164.380 116.300 164.640 ;
        RECT 116.360 164.380 116.620 164.640 ;
        RECT 116.680 164.380 116.940 164.640 ;
        RECT 117.000 164.380 117.260 164.640 ;
        RECT 117.320 164.380 117.580 164.640 ;
        RECT 85.610 163.870 85.870 164.130 ;
        RECT 89.290 163.870 89.550 164.130 ;
        RECT 95.730 163.870 95.990 164.130 ;
        RECT 94.350 163.530 94.610 163.790 ;
        RECT 75.490 162.850 75.750 163.110 ;
        RECT 76.870 162.850 77.130 163.110 ;
        RECT 79.170 162.850 79.430 163.110 ;
        RECT 111.830 163.530 112.090 163.790 ;
        RECT 108.150 162.850 108.410 163.110 ;
        RECT 82.850 162.170 83.110 162.430 ;
        RECT 84.230 162.170 84.490 162.430 ;
        RECT 93.890 162.170 94.150 162.430 ;
        RECT 109.530 162.170 109.790 162.430 ;
        RECT 115.050 162.170 115.310 162.430 ;
        RECT 76.515 161.660 76.775 161.920 ;
        RECT 76.835 161.660 77.095 161.920 ;
        RECT 77.155 161.660 77.415 161.920 ;
        RECT 77.475 161.660 77.735 161.920 ;
        RECT 77.795 161.660 78.055 161.920 ;
        RECT 88.590 161.660 88.850 161.920 ;
        RECT 88.910 161.660 89.170 161.920 ;
        RECT 89.230 161.660 89.490 161.920 ;
        RECT 89.550 161.660 89.810 161.920 ;
        RECT 89.870 161.660 90.130 161.920 ;
        RECT 100.665 161.660 100.925 161.920 ;
        RECT 100.985 161.660 101.245 161.920 ;
        RECT 101.305 161.660 101.565 161.920 ;
        RECT 101.625 161.660 101.885 161.920 ;
        RECT 101.945 161.660 102.205 161.920 ;
        RECT 112.740 161.660 113.000 161.920 ;
        RECT 113.060 161.660 113.320 161.920 ;
        RECT 113.380 161.660 113.640 161.920 ;
        RECT 113.700 161.660 113.960 161.920 ;
        RECT 114.020 161.660 114.280 161.920 ;
        RECT 84.230 161.150 84.490 161.410 ;
        RECT 106.310 161.150 106.570 161.410 ;
        RECT 114.590 161.150 114.850 161.410 ;
        RECT 102.630 160.810 102.890 161.070 ;
        RECT 115.050 160.470 115.310 160.730 ;
        RECT 102.170 160.130 102.430 160.390 ;
        RECT 103.090 160.130 103.350 160.390 ;
        RECT 108.610 160.130 108.870 160.390 ;
        RECT 109.530 160.130 109.790 160.390 ;
        RECT 110.450 160.130 110.710 160.390 ;
        RECT 87.910 159.450 88.170 159.710 ;
        RECT 103.550 159.450 103.810 159.710 ;
        RECT 79.815 158.940 80.075 159.200 ;
        RECT 80.135 158.940 80.395 159.200 ;
        RECT 80.455 158.940 80.715 159.200 ;
        RECT 80.775 158.940 81.035 159.200 ;
        RECT 81.095 158.940 81.355 159.200 ;
        RECT 91.890 158.940 92.150 159.200 ;
        RECT 92.210 158.940 92.470 159.200 ;
        RECT 92.530 158.940 92.790 159.200 ;
        RECT 92.850 158.940 93.110 159.200 ;
        RECT 93.170 158.940 93.430 159.200 ;
        RECT 103.965 158.940 104.225 159.200 ;
        RECT 104.285 158.940 104.545 159.200 ;
        RECT 104.605 158.940 104.865 159.200 ;
        RECT 104.925 158.940 105.185 159.200 ;
        RECT 105.245 158.940 105.505 159.200 ;
        RECT 116.040 158.940 116.300 159.200 ;
        RECT 116.360 158.940 116.620 159.200 ;
        RECT 116.680 158.940 116.940 159.200 ;
        RECT 117.000 158.940 117.260 159.200 ;
        RECT 117.320 158.940 117.580 159.200 ;
        RECT 102.170 158.430 102.430 158.690 ;
        RECT 82.850 158.090 83.110 158.350 ;
        RECT 95.730 158.090 95.990 158.350 ;
        RECT 82.390 157.750 82.650 158.010 ;
        RECT 85.610 157.410 85.870 157.670 ;
        RECT 93.430 157.750 93.690 158.010 ;
        RECT 103.090 157.750 103.350 158.010 ;
        RECT 87.910 157.410 88.170 157.670 ;
        RECT 79.170 156.730 79.430 156.990 ;
        RECT 90.210 157.070 90.470 157.330 ;
        RECT 102.630 157.070 102.890 157.330 ;
        RECT 104.930 157.410 105.190 157.670 ;
        RECT 109.530 157.750 109.790 158.010 ;
        RECT 115.050 157.750 115.310 158.010 ;
        RECT 118.730 157.750 118.990 158.010 ;
        RECT 108.610 157.410 108.870 157.670 ;
        RECT 110.910 157.410 111.170 157.670 ;
        RECT 115.510 157.410 115.770 157.670 ;
        RECT 94.350 156.730 94.610 156.990 ;
        RECT 103.090 156.730 103.350 156.990 ;
        RECT 104.470 156.730 104.730 156.990 ;
        RECT 110.450 156.730 110.710 156.990 ;
        RECT 76.515 156.220 76.775 156.480 ;
        RECT 76.835 156.220 77.095 156.480 ;
        RECT 77.155 156.220 77.415 156.480 ;
        RECT 77.475 156.220 77.735 156.480 ;
        RECT 77.795 156.220 78.055 156.480 ;
        RECT 88.590 156.220 88.850 156.480 ;
        RECT 88.910 156.220 89.170 156.480 ;
        RECT 89.230 156.220 89.490 156.480 ;
        RECT 89.550 156.220 89.810 156.480 ;
        RECT 89.870 156.220 90.130 156.480 ;
        RECT 100.665 156.220 100.925 156.480 ;
        RECT 100.985 156.220 101.245 156.480 ;
        RECT 101.305 156.220 101.565 156.480 ;
        RECT 101.625 156.220 101.885 156.480 ;
        RECT 101.945 156.220 102.205 156.480 ;
        RECT 112.740 156.220 113.000 156.480 ;
        RECT 113.060 156.220 113.320 156.480 ;
        RECT 113.380 156.220 113.640 156.480 ;
        RECT 113.700 156.220 113.960 156.480 ;
        RECT 114.020 156.220 114.280 156.480 ;
        RECT 15.245 147.590 15.980 148.210 ;
        RECT 20.425 149.845 20.685 150.105 ;
        RECT 19.630 147.565 19.960 147.865 ;
        RECT 82.390 155.710 82.650 155.970 ;
        RECT 94.350 155.710 94.610 155.970 ;
        RECT 103.090 155.710 103.350 155.970 ;
        RECT 104.470 155.710 104.730 155.970 ;
        RECT 108.610 155.710 108.870 155.970 ;
        RECT 115.510 155.710 115.770 155.970 ;
        RECT 117.810 155.710 118.070 155.970 ;
        RECT 106.770 155.370 107.030 155.630 ;
        RECT 75.490 155.030 75.750 155.290 ;
        RECT 93.890 155.030 94.150 155.290 ;
        RECT 75.030 154.350 75.290 154.610 ;
        RECT 82.850 154.690 83.110 154.950 ;
        RECT 84.230 154.690 84.490 154.950 ;
        RECT 84.690 154.010 84.950 154.270 ;
        RECT 95.730 154.350 95.990 154.610 ;
        RECT 108.150 155.030 108.410 155.290 ;
        RECT 93.890 154.010 94.150 154.270 ;
        RECT 109.530 154.690 109.790 154.950 ;
        RECT 103.550 154.350 103.810 154.610 ;
        RECT 102.170 154.010 102.430 154.270 ;
        RECT 103.090 154.010 103.350 154.270 ;
        RECT 115.050 154.350 115.310 154.610 ;
        RECT 79.815 153.500 80.075 153.760 ;
        RECT 80.135 153.500 80.395 153.760 ;
        RECT 80.455 153.500 80.715 153.760 ;
        RECT 80.775 153.500 81.035 153.760 ;
        RECT 81.095 153.500 81.355 153.760 ;
        RECT 91.890 153.500 92.150 153.760 ;
        RECT 92.210 153.500 92.470 153.760 ;
        RECT 92.530 153.500 92.790 153.760 ;
        RECT 92.850 153.500 93.110 153.760 ;
        RECT 93.170 153.500 93.430 153.760 ;
        RECT 103.965 153.500 104.225 153.760 ;
        RECT 104.285 153.500 104.545 153.760 ;
        RECT 104.605 153.500 104.865 153.760 ;
        RECT 104.925 153.500 105.185 153.760 ;
        RECT 105.245 153.500 105.505 153.760 ;
        RECT 116.040 153.500 116.300 153.760 ;
        RECT 116.360 153.500 116.620 153.760 ;
        RECT 116.680 153.500 116.940 153.760 ;
        RECT 117.000 153.500 117.260 153.760 ;
        RECT 117.320 153.500 117.580 153.760 ;
        RECT 75.030 152.990 75.290 153.250 ;
        RECT 84.690 152.990 84.950 153.250 ;
        RECT 96.650 152.650 96.910 152.910 ;
        RECT 107.230 152.990 107.490 153.250 ;
        RECT 110.910 152.990 111.170 153.250 ;
        RECT 115.050 152.990 115.310 153.250 ;
        RECT 119.190 152.990 119.450 153.250 ;
        RECT 120.110 152.990 120.370 153.250 ;
        RECT 102.170 152.650 102.430 152.910 ;
        RECT 81.470 151.970 81.730 152.230 ;
        RECT 93.890 151.970 94.150 152.230 ;
        RECT 82.850 151.630 83.110 151.890 ;
        RECT 86.070 151.630 86.330 151.890 ;
        RECT 84.230 151.290 84.490 151.550 ;
        RECT 103.090 152.310 103.350 152.570 ;
        RECT 105.390 152.310 105.650 152.570 ;
        RECT 102.630 151.630 102.890 151.890 ;
        RECT 114.590 151.290 114.850 151.550 ;
        RECT 76.515 150.780 76.775 151.040 ;
        RECT 76.835 150.780 77.095 151.040 ;
        RECT 77.155 150.780 77.415 151.040 ;
        RECT 77.475 150.780 77.735 151.040 ;
        RECT 77.795 150.780 78.055 151.040 ;
        RECT 88.590 150.780 88.850 151.040 ;
        RECT 88.910 150.780 89.170 151.040 ;
        RECT 89.230 150.780 89.490 151.040 ;
        RECT 89.550 150.780 89.810 151.040 ;
        RECT 89.870 150.780 90.130 151.040 ;
        RECT 100.665 150.780 100.925 151.040 ;
        RECT 100.985 150.780 101.245 151.040 ;
        RECT 101.305 150.780 101.565 151.040 ;
        RECT 101.625 150.780 101.885 151.040 ;
        RECT 101.945 150.780 102.205 151.040 ;
        RECT 112.740 150.780 113.000 151.040 ;
        RECT 113.060 150.780 113.320 151.040 ;
        RECT 113.380 150.780 113.640 151.040 ;
        RECT 113.700 150.780 113.960 151.040 ;
        RECT 114.020 150.780 114.280 151.040 ;
        RECT 81.930 150.270 82.190 150.530 ;
        RECT 93.890 150.270 94.150 150.530 ;
        RECT 102.630 150.270 102.890 150.530 ;
        RECT 105.390 150.270 105.650 150.530 ;
        RECT 114.590 150.270 114.850 150.530 ;
        RECT 84.230 149.590 84.490 149.850 ;
        RECT 107.230 149.930 107.490 150.190 ;
        RECT 81.930 149.250 82.190 149.510 ;
        RECT 85.610 148.910 85.870 149.170 ;
        RECT 87.450 148.910 87.710 149.170 ;
        RECT 106.770 149.250 107.030 149.510 ;
        RECT 110.910 149.590 111.170 149.850 ;
        RECT 117.810 149.590 118.070 149.850 ;
        RECT 109.530 148.910 109.790 149.170 ;
        RECT 109.070 148.570 109.330 148.830 ;
        RECT 49.415 147.950 49.895 148.430 ;
        RECT 79.815 148.060 80.075 148.320 ;
        RECT 80.135 148.060 80.395 148.320 ;
        RECT 80.455 148.060 80.715 148.320 ;
        RECT 80.775 148.060 81.035 148.320 ;
        RECT 81.095 148.060 81.355 148.320 ;
        RECT 91.890 148.060 92.150 148.320 ;
        RECT 92.210 148.060 92.470 148.320 ;
        RECT 92.530 148.060 92.790 148.320 ;
        RECT 92.850 148.060 93.110 148.320 ;
        RECT 93.170 148.060 93.430 148.320 ;
        RECT 103.965 148.060 104.225 148.320 ;
        RECT 104.285 148.060 104.545 148.320 ;
        RECT 104.605 148.060 104.865 148.320 ;
        RECT 104.925 148.060 105.185 148.320 ;
        RECT 105.245 148.060 105.505 148.320 ;
        RECT 116.040 148.060 116.300 148.320 ;
        RECT 116.360 148.060 116.620 148.320 ;
        RECT 116.680 148.060 116.940 148.320 ;
        RECT 117.000 148.060 117.260 148.320 ;
        RECT 117.320 148.060 117.580 148.320 ;
        RECT 21.090 143.000 21.350 143.260 ;
        RECT 19.840 140.425 20.120 140.705 ;
        RECT 18.915 139.155 19.175 139.415 ;
        RECT 25.545 143.440 26.260 144.195 ;
        RECT 21.350 135.295 21.610 135.555 ;
        RECT 24.500 135.385 24.780 135.665 ;
        RECT 21.980 133.855 22.310 134.135 ;
        RECT 24.040 133.875 24.300 134.135 ;
        RECT 17.640 131.180 17.900 131.440 ;
        RECT 19.640 131.075 19.900 131.335 ;
        RECT 23.960 130.465 24.250 130.735 ;
        RECT 13.070 123.935 13.935 124.915 ;
        RECT 14.650 109.065 15.280 109.635 ;
        RECT 20.205 111.875 20.465 112.135 ;
        RECT 19.410 109.595 19.740 109.895 ;
        RECT 20.870 105.030 21.130 105.290 ;
        RECT 19.620 102.455 19.900 102.735 ;
        RECT 18.695 101.185 18.955 101.445 ;
        RECT 25.325 105.470 26.040 106.225 ;
        RECT 21.130 97.325 21.390 97.585 ;
        RECT 24.280 97.415 24.560 97.695 ;
        RECT 21.760 95.885 22.090 96.165 ;
        RECT 23.820 95.905 24.080 96.165 ;
        RECT 19.420 93.105 19.680 93.365 ;
        RECT 23.740 92.495 24.030 92.765 ;
        RECT 1.365 82.730 2.055 83.240 ;
        RECT 49.350 88.610 50.010 89.310 ;
        RECT 101.235 88.810 101.495 89.070 ;
        RECT 101.555 88.810 101.815 89.070 ;
        RECT 101.875 88.810 102.135 89.070 ;
        RECT 102.195 88.810 102.455 89.070 ;
        RECT 102.515 88.810 102.775 89.070 ;
        RECT 116.530 88.810 116.790 89.070 ;
        RECT 116.850 88.810 117.110 89.070 ;
        RECT 117.170 88.810 117.430 89.070 ;
        RECT 117.490 88.810 117.750 89.070 ;
        RECT 117.810 88.810 118.070 89.070 ;
        RECT 131.825 88.810 132.085 89.070 ;
        RECT 132.145 88.810 132.405 89.070 ;
        RECT 132.465 88.810 132.725 89.070 ;
        RECT 132.785 88.810 133.045 89.070 ;
        RECT 133.105 88.810 133.365 89.070 ;
        RECT 147.120 88.810 147.380 89.070 ;
        RECT 147.440 88.810 147.700 89.070 ;
        RECT 147.760 88.810 148.020 89.070 ;
        RECT 148.080 88.810 148.340 89.070 ;
        RECT 148.400 88.810 148.660 89.070 ;
        RECT 103.580 88.300 103.840 88.560 ;
        RECT 139.460 88.300 139.720 88.560 ;
        RECT 151.880 87.960 152.140 88.220 ;
        RECT 106.340 87.620 106.600 87.880 ;
        RECT 140.380 87.620 140.640 87.880 ;
        RECT 145.900 86.940 146.160 87.200 ;
        RECT 97.935 86.090 98.195 86.350 ;
        RECT 98.255 86.090 98.515 86.350 ;
        RECT 98.575 86.090 98.835 86.350 ;
        RECT 98.895 86.090 99.155 86.350 ;
        RECT 99.215 86.090 99.475 86.350 ;
        RECT 113.230 86.090 113.490 86.350 ;
        RECT 113.550 86.090 113.810 86.350 ;
        RECT 113.870 86.090 114.130 86.350 ;
        RECT 114.190 86.090 114.450 86.350 ;
        RECT 114.510 86.090 114.770 86.350 ;
        RECT 128.525 86.090 128.785 86.350 ;
        RECT 128.845 86.090 129.105 86.350 ;
        RECT 129.165 86.090 129.425 86.350 ;
        RECT 129.485 86.090 129.745 86.350 ;
        RECT 129.805 86.090 130.065 86.350 ;
        RECT 143.820 86.090 144.080 86.350 ;
        RECT 144.140 86.090 144.400 86.350 ;
        RECT 144.460 86.090 144.720 86.350 ;
        RECT 144.780 86.090 145.040 86.350 ;
        RECT 145.100 86.090 145.360 86.350 ;
        RECT 118.300 84.900 118.560 85.160 ;
        RECT 125.660 84.900 125.920 85.160 ;
        RECT 121.980 84.560 122.240 84.820 ;
        RECT 122.440 84.560 122.700 84.820 ;
        RECT 126.120 84.560 126.380 84.820 ;
        RECT 122.900 83.880 123.160 84.140 ;
        RECT 124.740 83.880 125.000 84.140 ;
        RECT 127.500 83.880 127.760 84.140 ;
        RECT 143.600 84.560 143.860 84.820 ;
        RECT 145.440 83.880 145.700 84.140 ;
        RECT 101.235 83.370 101.495 83.630 ;
        RECT 101.555 83.370 101.815 83.630 ;
        RECT 101.875 83.370 102.135 83.630 ;
        RECT 102.195 83.370 102.455 83.630 ;
        RECT 102.515 83.370 102.775 83.630 ;
        RECT 116.530 83.370 116.790 83.630 ;
        RECT 116.850 83.370 117.110 83.630 ;
        RECT 117.170 83.370 117.430 83.630 ;
        RECT 117.490 83.370 117.750 83.630 ;
        RECT 117.810 83.370 118.070 83.630 ;
        RECT 131.825 83.370 132.085 83.630 ;
        RECT 132.145 83.370 132.405 83.630 ;
        RECT 132.465 83.370 132.725 83.630 ;
        RECT 132.785 83.370 133.045 83.630 ;
        RECT 133.105 83.370 133.365 83.630 ;
        RECT 147.120 83.370 147.380 83.630 ;
        RECT 147.440 83.370 147.700 83.630 ;
        RECT 147.760 83.370 148.020 83.630 ;
        RECT 148.080 83.370 148.340 83.630 ;
        RECT 148.400 83.370 148.660 83.630 ;
        RECT 122.440 82.860 122.700 83.120 ;
        RECT 118.760 82.520 119.020 82.780 ;
        RECT 113.240 81.840 113.500 82.100 ;
        RECT 115.080 81.840 115.340 82.100 ;
        RECT 118.300 81.840 118.560 82.100 ;
        RECT 121.980 82.520 122.240 82.780 ;
        RECT 125.660 82.520 125.920 82.780 ;
        RECT 127.960 82.520 128.220 82.780 ;
        RECT 124.740 81.840 125.000 82.100 ;
        RECT 143.600 82.860 143.860 83.120 ;
        RECT 133.940 82.180 134.200 82.440 ;
        RECT 142.680 82.180 142.940 82.440 ;
        RECT 145.900 82.180 146.160 82.440 ;
        RECT 136.240 81.840 136.500 82.100 ;
        RECT 134.860 81.500 135.120 81.760 ;
        RECT 115.540 81.160 115.800 81.420 ;
        RECT 121.520 81.160 121.780 81.420 ;
        RECT 122.440 81.160 122.700 81.420 ;
        RECT 137.160 81.160 137.420 81.420 ;
        RECT 97.935 80.650 98.195 80.910 ;
        RECT 98.255 80.650 98.515 80.910 ;
        RECT 98.575 80.650 98.835 80.910 ;
        RECT 98.895 80.650 99.155 80.910 ;
        RECT 99.215 80.650 99.475 80.910 ;
        RECT 113.230 80.650 113.490 80.910 ;
        RECT 113.550 80.650 113.810 80.910 ;
        RECT 113.870 80.650 114.130 80.910 ;
        RECT 114.190 80.650 114.450 80.910 ;
        RECT 114.510 80.650 114.770 80.910 ;
        RECT 128.525 80.650 128.785 80.910 ;
        RECT 128.845 80.650 129.105 80.910 ;
        RECT 129.165 80.650 129.425 80.910 ;
        RECT 129.485 80.650 129.745 80.910 ;
        RECT 129.805 80.650 130.065 80.910 ;
        RECT 143.820 80.650 144.080 80.910 ;
        RECT 144.140 80.650 144.400 80.910 ;
        RECT 144.460 80.650 144.720 80.910 ;
        RECT 144.780 80.650 145.040 80.910 ;
        RECT 145.100 80.650 145.360 80.910 ;
        RECT 122.900 80.140 123.160 80.400 ;
        RECT 110.940 79.460 111.200 79.720 ;
        RECT 118.300 79.460 118.560 79.720 ;
        RECT 115.080 78.780 115.340 79.040 ;
        RECT 119.220 79.120 119.480 79.380 ;
        RECT 127.960 80.140 128.220 80.400 ;
        RECT 133.940 80.140 134.200 80.400 ;
        RECT 127.500 79.800 127.760 80.060 ;
        RECT 137.620 80.140 137.880 80.400 ;
        RECT 145.440 80.140 145.700 80.400 ;
        RECT 124.280 79.120 124.540 79.380 ;
        RECT 122.440 78.780 122.700 79.040 ;
        RECT 126.120 78.780 126.380 79.040 ;
        RECT 127.500 78.780 127.760 79.040 ;
        RECT 131.180 79.120 131.440 79.380 ;
        RECT 130.720 78.780 130.980 79.040 ;
        RECT 134.860 79.120 135.120 79.380 ;
        RECT 136.240 79.120 136.500 79.380 ;
        RECT 115.540 78.440 115.800 78.700 ;
        RECT 121.060 78.440 121.320 78.700 ;
        RECT 133.710 78.440 133.970 78.700 ;
        RECT 135.320 78.440 135.580 78.700 ;
        RECT 145.900 79.120 146.160 79.380 ;
        RECT 137.160 78.440 137.420 78.700 ;
        RECT 143.140 78.440 143.400 78.700 ;
        RECT 101.235 77.930 101.495 78.190 ;
        RECT 101.555 77.930 101.815 78.190 ;
        RECT 101.875 77.930 102.135 78.190 ;
        RECT 102.195 77.930 102.455 78.190 ;
        RECT 102.515 77.930 102.775 78.190 ;
        RECT 116.530 77.930 116.790 78.190 ;
        RECT 116.850 77.930 117.110 78.190 ;
        RECT 117.170 77.930 117.430 78.190 ;
        RECT 117.490 77.930 117.750 78.190 ;
        RECT 117.810 77.930 118.070 78.190 ;
        RECT 131.825 77.930 132.085 78.190 ;
        RECT 132.145 77.930 132.405 78.190 ;
        RECT 132.465 77.930 132.725 78.190 ;
        RECT 132.785 77.930 133.045 78.190 ;
        RECT 133.105 77.930 133.365 78.190 ;
        RECT 147.120 77.930 147.380 78.190 ;
        RECT 147.440 77.930 147.700 78.190 ;
        RECT 147.760 77.930 148.020 78.190 ;
        RECT 148.080 77.930 148.340 78.190 ;
        RECT 148.400 77.930 148.660 78.190 ;
        RECT 7.575 72.720 7.985 73.025 ;
        RECT 23.500 71.940 23.760 72.200 ;
        RECT 32.960 71.970 33.340 72.280 ;
        RECT 7.640 68.595 7.935 68.975 ;
        RECT 27.570 69.705 27.905 70.030 ;
        RECT 27.470 67.450 27.770 67.740 ;
        RECT 115.080 76.740 115.340 77.000 ;
        RECT 118.300 76.740 118.560 77.000 ;
        RECT 121.520 77.420 121.780 77.680 ;
        RECT 121.980 77.420 122.240 77.680 ;
        RECT 133.020 77.420 133.280 77.680 ;
        RECT 121.060 76.740 121.320 77.000 ;
        RECT 135.780 77.420 136.040 77.680 ;
        RECT 136.700 77.420 136.960 77.680 ;
        RECT 113.240 76.400 113.500 76.660 ;
        RECT 127.500 76.400 127.760 76.660 ;
        RECT 131.180 76.400 131.440 76.660 ;
        RECT 133.480 76.740 133.740 77.000 ;
        RECT 135.320 76.740 135.580 77.000 ;
        RECT 136.240 76.740 136.500 77.000 ;
        RECT 137.620 76.740 137.880 77.000 ;
        RECT 140.380 76.740 140.640 77.000 ;
        RECT 145.440 77.420 145.700 77.680 ;
        RECT 107.260 75.720 107.520 75.980 ;
        RECT 121.520 75.720 121.780 75.980 ;
        RECT 127.040 75.720 127.300 75.980 ;
        RECT 143.140 76.400 143.400 76.660 ;
        RECT 139.000 75.720 139.260 75.980 ;
        RECT 141.300 75.720 141.560 75.980 ;
        RECT 141.760 75.720 142.020 75.980 ;
        RECT 142.680 75.720 142.940 75.980 ;
        RECT 145.440 75.720 145.700 75.980 ;
        RECT 146.820 75.720 147.080 75.980 ;
        RECT 97.935 75.210 98.195 75.470 ;
        RECT 98.255 75.210 98.515 75.470 ;
        RECT 98.575 75.210 98.835 75.470 ;
        RECT 98.895 75.210 99.155 75.470 ;
        RECT 99.215 75.210 99.475 75.470 ;
        RECT 113.230 75.210 113.490 75.470 ;
        RECT 113.550 75.210 113.810 75.470 ;
        RECT 113.870 75.210 114.130 75.470 ;
        RECT 114.190 75.210 114.450 75.470 ;
        RECT 114.510 75.210 114.770 75.470 ;
        RECT 128.525 75.210 128.785 75.470 ;
        RECT 128.845 75.210 129.105 75.470 ;
        RECT 129.165 75.210 129.425 75.470 ;
        RECT 129.485 75.210 129.745 75.470 ;
        RECT 129.805 75.210 130.065 75.470 ;
        RECT 143.820 75.210 144.080 75.470 ;
        RECT 144.140 75.210 144.400 75.470 ;
        RECT 144.460 75.210 144.720 75.470 ;
        RECT 144.780 75.210 145.040 75.470 ;
        RECT 145.100 75.210 145.360 75.470 ;
        RECT 105.880 74.700 106.140 74.960 ;
        RECT 115.540 74.700 115.800 74.960 ;
        RECT 118.760 74.700 119.020 74.960 ;
        RECT 130.720 74.700 130.980 74.960 ;
        RECT 139.000 74.700 139.260 74.960 ;
        RECT 141.300 74.700 141.560 74.960 ;
        RECT 146.820 74.700 147.080 74.960 ;
        RECT 119.220 74.360 119.480 74.620 ;
        RECT 118.300 74.020 118.560 74.280 ;
        RECT 135.780 74.360 136.040 74.620 ;
        RECT 110.940 73.680 111.200 73.940 ;
        RECT 107.260 73.340 107.520 73.600 ;
        RECT 109.100 73.340 109.360 73.600 ;
        RECT 120.600 73.680 120.860 73.940 ;
        RECT 121.520 73.680 121.780 73.940 ;
        RECT 121.980 73.680 122.240 73.940 ;
        RECT 122.440 73.680 122.700 73.940 ;
        RECT 138.080 74.020 138.340 74.280 ;
        RECT 127.040 73.340 127.300 73.600 ;
        RECT 127.500 73.340 127.760 73.600 ;
        RECT 137.620 73.680 137.880 73.940 ;
        RECT 141.300 73.680 141.560 73.940 ;
        RECT 142.680 74.360 142.940 74.620 ;
        RECT 142.220 73.680 142.480 73.940 ;
        RECT 143.140 73.680 143.400 73.940 ;
        RECT 143.600 73.680 143.860 73.940 ;
        RECT 118.760 73.000 119.020 73.260 ;
        RECT 133.480 73.340 133.740 73.600 ;
        RECT 135.320 73.000 135.580 73.260 ;
        RECT 145.900 73.680 146.160 73.940 ;
        RECT 146.360 73.680 146.620 73.940 ;
        RECT 140.840 73.000 141.100 73.260 ;
        RECT 143.140 73.000 143.400 73.260 ;
        RECT 145.900 73.000 146.160 73.260 ;
        RECT 101.235 72.490 101.495 72.750 ;
        RECT 101.555 72.490 101.815 72.750 ;
        RECT 101.875 72.490 102.135 72.750 ;
        RECT 102.195 72.490 102.455 72.750 ;
        RECT 102.515 72.490 102.775 72.750 ;
        RECT 116.530 72.490 116.790 72.750 ;
        RECT 116.850 72.490 117.110 72.750 ;
        RECT 117.170 72.490 117.430 72.750 ;
        RECT 117.490 72.490 117.750 72.750 ;
        RECT 117.810 72.490 118.070 72.750 ;
        RECT 131.825 72.490 132.085 72.750 ;
        RECT 132.145 72.490 132.405 72.750 ;
        RECT 132.465 72.490 132.725 72.750 ;
        RECT 132.785 72.490 133.045 72.750 ;
        RECT 133.105 72.490 133.365 72.750 ;
        RECT 147.120 72.490 147.380 72.750 ;
        RECT 147.440 72.490 147.700 72.750 ;
        RECT 147.760 72.490 148.020 72.750 ;
        RECT 148.080 72.490 148.340 72.750 ;
        RECT 148.400 72.490 148.660 72.750 ;
        RECT 109.100 71.980 109.360 72.240 ;
        RECT 115.080 71.980 115.340 72.240 ;
        RECT 109.560 71.300 109.820 71.560 ;
        RECT 112.780 71.300 113.040 71.560 ;
        RECT 118.760 71.640 119.020 71.900 ;
        RECT 115.080 70.280 115.340 70.540 ;
        RECT 120.600 71.300 120.860 71.560 ;
        RECT 127.500 71.640 127.760 71.900 ;
        RECT 127.040 71.300 127.300 71.560 ;
        RECT 136.700 71.980 136.960 72.240 ;
        RECT 139.000 71.980 139.260 72.240 ;
        RECT 140.380 71.980 140.640 72.240 ;
        RECT 145.440 71.980 145.700 72.240 ;
        RECT 134.400 71.300 134.660 71.560 ;
        RECT 148.660 71.640 148.920 71.900 ;
        RECT 118.300 70.960 118.560 71.220 ;
        RECT 122.440 70.960 122.700 71.220 ;
        RECT 137.620 71.300 137.880 71.560 ;
        RECT 119.220 70.620 119.480 70.880 ;
        RECT 138.540 70.620 138.800 70.880 ;
        RECT 140.380 70.960 140.640 71.220 ;
        RECT 140.840 70.620 141.100 70.880 ;
        RECT 143.140 71.300 143.400 71.560 ;
        RECT 145.900 71.300 146.160 71.560 ;
        RECT 146.820 71.300 147.080 71.560 ;
        RECT 147.280 71.300 147.540 71.560 ;
        RECT 142.680 70.960 142.940 71.220 ;
        RECT 143.600 70.960 143.860 71.220 ;
        RECT 127.500 70.280 127.760 70.540 ;
        RECT 133.480 70.280 133.740 70.540 ;
        RECT 140.380 70.280 140.640 70.540 ;
        RECT 143.140 70.620 143.400 70.880 ;
        RECT 150.500 70.960 150.760 71.220 ;
        RECT 145.440 70.280 145.700 70.540 ;
        RECT 97.935 69.770 98.195 70.030 ;
        RECT 98.255 69.770 98.515 70.030 ;
        RECT 98.575 69.770 98.835 70.030 ;
        RECT 98.895 69.770 99.155 70.030 ;
        RECT 99.215 69.770 99.475 70.030 ;
        RECT 113.230 69.770 113.490 70.030 ;
        RECT 113.550 69.770 113.810 70.030 ;
        RECT 113.870 69.770 114.130 70.030 ;
        RECT 114.190 69.770 114.450 70.030 ;
        RECT 114.510 69.770 114.770 70.030 ;
        RECT 128.525 69.770 128.785 70.030 ;
        RECT 128.845 69.770 129.105 70.030 ;
        RECT 129.165 69.770 129.425 70.030 ;
        RECT 129.485 69.770 129.745 70.030 ;
        RECT 129.805 69.770 130.065 70.030 ;
        RECT 143.820 69.770 144.080 70.030 ;
        RECT 144.140 69.770 144.400 70.030 ;
        RECT 144.460 69.770 144.720 70.030 ;
        RECT 144.780 69.770 145.040 70.030 ;
        RECT 145.100 69.770 145.360 70.030 ;
        RECT 118.300 69.260 118.560 69.520 ;
        RECT 134.400 69.260 134.660 69.520 ;
        RECT 135.320 69.260 135.580 69.520 ;
        RECT 138.080 69.260 138.340 69.520 ;
        RECT 138.540 69.260 138.800 69.520 ;
        RECT 140.380 69.260 140.640 69.520 ;
        RECT 144.060 69.260 144.320 69.520 ;
        RECT 146.360 69.260 146.620 69.520 ;
        RECT 137.620 68.920 137.880 69.180 ;
        RECT 110.940 68.580 111.200 68.840 ;
        RECT 115.080 68.580 115.340 68.840 ;
        RECT 103.580 68.240 103.840 68.500 ;
        RECT 115.080 67.900 115.340 68.160 ;
        RECT 122.440 68.240 122.700 68.500 ;
        RECT 140.840 68.580 141.100 68.840 ;
        RECT 143.600 68.580 143.860 68.840 ;
        RECT 145.440 68.580 145.700 68.840 ;
        RECT 100.360 67.560 100.620 67.820 ;
        RECT 121.060 67.560 121.320 67.820 ;
        RECT 135.320 67.560 135.580 67.820 ;
        RECT 141.760 68.240 142.020 68.500 ;
        RECT 143.140 68.240 143.400 68.500 ;
        RECT 148.660 68.240 148.920 68.500 ;
        RECT 142.680 67.560 142.940 67.820 ;
        RECT 144.980 67.560 145.240 67.820 ;
        RECT 145.440 67.560 145.700 67.820 ;
        RECT 145.900 67.560 146.160 67.820 ;
        RECT 147.280 67.560 147.540 67.820 ;
        RECT 101.235 67.050 101.495 67.310 ;
        RECT 101.555 67.050 101.815 67.310 ;
        RECT 101.875 67.050 102.135 67.310 ;
        RECT 102.195 67.050 102.455 67.310 ;
        RECT 102.515 67.050 102.775 67.310 ;
        RECT 116.530 67.050 116.790 67.310 ;
        RECT 116.850 67.050 117.110 67.310 ;
        RECT 117.170 67.050 117.430 67.310 ;
        RECT 117.490 67.050 117.750 67.310 ;
        RECT 117.810 67.050 118.070 67.310 ;
        RECT 131.825 67.050 132.085 67.310 ;
        RECT 132.145 67.050 132.405 67.310 ;
        RECT 132.465 67.050 132.725 67.310 ;
        RECT 132.785 67.050 133.045 67.310 ;
        RECT 133.105 67.050 133.365 67.310 ;
        RECT 147.120 67.050 147.380 67.310 ;
        RECT 147.440 67.050 147.700 67.310 ;
        RECT 147.760 67.050 148.020 67.310 ;
        RECT 148.080 67.050 148.340 67.310 ;
        RECT 148.400 67.050 148.660 67.310 ;
        RECT 35.225 65.665 35.495 65.925 ;
        RECT 34.540 64.690 34.850 64.970 ;
        RECT 19.080 63.390 19.420 63.660 ;
        RECT 7.395 57.315 8.255 58.175 ;
        RECT 23.180 56.600 23.630 57.180 ;
        RECT 27.730 63.340 28.065 63.665 ;
        RECT 53.395 61.225 53.760 61.605 ;
        RECT 28.780 59.195 29.190 59.545 ;
        RECT 34.220 59.225 34.670 59.575 ;
        RECT 26.535 57.930 26.900 58.460 ;
        RECT 109.560 66.540 109.820 66.800 ;
        RECT 100.360 66.200 100.620 66.460 ;
        RECT 115.080 66.540 115.340 66.800 ;
        RECT 122.440 66.540 122.700 66.800 ;
        RECT 127.960 66.200 128.220 66.460 ;
        RECT 101.740 64.840 102.000 65.100 ;
        RECT 103.120 64.840 103.380 65.100 ;
        RECT 124.280 65.860 124.540 66.120 ;
        RECT 138.080 66.540 138.340 66.800 ;
        RECT 143.140 66.540 143.400 66.800 ;
        RECT 134.400 65.860 134.660 66.120 ;
        RECT 127.500 65.520 127.760 65.780 ;
        RECT 139.920 65.860 140.180 66.120 ;
        RECT 144.060 65.860 144.320 66.120 ;
        RECT 145.440 65.860 145.700 66.120 ;
        RECT 145.900 65.860 146.160 66.120 ;
        RECT 135.320 65.520 135.580 65.780 ;
        RECT 142.220 65.520 142.480 65.780 ;
        RECT 141.300 65.180 141.560 65.440 ;
        RECT 107.260 64.840 107.520 65.100 ;
        RECT 122.440 64.840 122.700 65.100 ;
        RECT 138.080 64.840 138.340 65.100 ;
        RECT 140.840 64.840 141.100 65.100 ;
        RECT 142.680 64.840 142.940 65.100 ;
        RECT 143.140 64.840 143.400 65.100 ;
        RECT 144.060 64.840 144.320 65.100 ;
        RECT 150.960 64.840 151.220 65.100 ;
        RECT 97.935 64.330 98.195 64.590 ;
        RECT 98.255 64.330 98.515 64.590 ;
        RECT 98.575 64.330 98.835 64.590 ;
        RECT 98.895 64.330 99.155 64.590 ;
        RECT 99.215 64.330 99.475 64.590 ;
        RECT 113.230 64.330 113.490 64.590 ;
        RECT 113.550 64.330 113.810 64.590 ;
        RECT 113.870 64.330 114.130 64.590 ;
        RECT 114.190 64.330 114.450 64.590 ;
        RECT 114.510 64.330 114.770 64.590 ;
        RECT 128.525 64.330 128.785 64.590 ;
        RECT 128.845 64.330 129.105 64.590 ;
        RECT 129.165 64.330 129.425 64.590 ;
        RECT 129.485 64.330 129.745 64.590 ;
        RECT 129.805 64.330 130.065 64.590 ;
        RECT 143.820 64.330 144.080 64.590 ;
        RECT 144.140 64.330 144.400 64.590 ;
        RECT 144.460 64.330 144.720 64.590 ;
        RECT 144.780 64.330 145.040 64.590 ;
        RECT 145.100 64.330 145.360 64.590 ;
        RECT 101.740 63.820 102.000 64.080 ;
        RECT 110.940 63.820 111.200 64.080 ;
        RECT 122.440 63.820 122.700 64.080 ;
        RECT 127.960 63.820 128.220 64.080 ;
        RECT 146.360 63.820 146.620 64.080 ;
        RECT 107.260 63.140 107.520 63.400 ;
        RECT 93.000 62.120 93.260 62.380 ;
        RECT 100.360 62.460 100.620 62.720 ;
        RECT 112.780 62.800 113.040 63.060 ;
        RECT 121.060 63.140 121.320 63.400 ;
        RECT 143.140 63.480 143.400 63.740 ;
        RECT 103.120 62.120 103.380 62.380 ;
        RECT 105.880 62.120 106.140 62.380 ;
        RECT 107.260 62.120 107.520 62.380 ;
        RECT 107.720 62.120 107.980 62.380 ;
        RECT 113.700 62.460 113.960 62.720 ;
        RECT 114.160 62.460 114.420 62.720 ;
        RECT 146.360 62.800 146.620 63.060 ;
        RECT 121.980 62.120 122.240 62.380 ;
        RECT 126.120 62.120 126.380 62.380 ;
        RECT 142.680 62.120 142.940 62.380 ;
        RECT 101.235 61.610 101.495 61.870 ;
        RECT 101.555 61.610 101.815 61.870 ;
        RECT 101.875 61.610 102.135 61.870 ;
        RECT 102.195 61.610 102.455 61.870 ;
        RECT 102.515 61.610 102.775 61.870 ;
        RECT 116.530 61.610 116.790 61.870 ;
        RECT 116.850 61.610 117.110 61.870 ;
        RECT 117.170 61.610 117.430 61.870 ;
        RECT 117.490 61.610 117.750 61.870 ;
        RECT 117.810 61.610 118.070 61.870 ;
        RECT 131.825 61.610 132.085 61.870 ;
        RECT 132.145 61.610 132.405 61.870 ;
        RECT 132.465 61.610 132.725 61.870 ;
        RECT 132.785 61.610 133.045 61.870 ;
        RECT 133.105 61.610 133.365 61.870 ;
        RECT 147.120 61.610 147.380 61.870 ;
        RECT 147.440 61.610 147.700 61.870 ;
        RECT 147.760 61.610 148.020 61.870 ;
        RECT 148.080 61.610 148.340 61.870 ;
        RECT 148.400 61.610 148.660 61.870 ;
        RECT 55.655 56.860 56.090 57.345 ;
        RECT 93.000 61.100 93.260 61.360 ;
        RECT 95.760 61.100 96.020 61.360 ;
        RECT 100.360 61.100 100.620 61.360 ;
        RECT 103.580 61.100 103.840 61.360 ;
        RECT 107.260 61.100 107.520 61.360 ;
        RECT 114.160 61.100 114.420 61.360 ;
        RECT 121.980 61.100 122.240 61.360 ;
        RECT 138.080 61.100 138.340 61.360 ;
        RECT 146.360 61.100 146.620 61.360 ;
        RECT 98.060 60.420 98.320 60.680 ;
        RECT 99.440 60.420 99.700 60.680 ;
        RECT 99.900 60.420 100.160 60.680 ;
        RECT 102.200 60.420 102.460 60.680 ;
        RECT 104.960 60.420 105.220 60.680 ;
        RECT 106.800 60.420 107.060 60.680 ;
        RECT 107.260 60.420 107.520 60.680 ;
        RECT 115.540 60.760 115.800 61.020 ;
        RECT 100.820 60.080 101.080 60.340 ;
        RECT 113.700 60.420 113.960 60.680 ;
        RECT 127.040 60.420 127.300 60.680 ;
        RECT 145.900 60.420 146.160 60.680 ;
        RECT 150.040 60.080 150.300 60.340 ;
        RECT 105.880 59.740 106.140 60.000 ;
        RECT 96.680 59.400 96.940 59.660 ;
        RECT 99.440 59.400 99.700 59.660 ;
        RECT 108.640 59.400 108.900 59.660 ;
        RECT 123.820 59.400 124.080 59.660 ;
        RECT 147.740 59.400 148.000 59.660 ;
        RECT 97.935 58.890 98.195 59.150 ;
        RECT 98.255 58.890 98.515 59.150 ;
        RECT 98.575 58.890 98.835 59.150 ;
        RECT 98.895 58.890 99.155 59.150 ;
        RECT 99.215 58.890 99.475 59.150 ;
        RECT 113.230 58.890 113.490 59.150 ;
        RECT 113.550 58.890 113.810 59.150 ;
        RECT 113.870 58.890 114.130 59.150 ;
        RECT 114.190 58.890 114.450 59.150 ;
        RECT 114.510 58.890 114.770 59.150 ;
        RECT 128.525 58.890 128.785 59.150 ;
        RECT 128.845 58.890 129.105 59.150 ;
        RECT 129.165 58.890 129.425 59.150 ;
        RECT 129.485 58.890 129.745 59.150 ;
        RECT 129.805 58.890 130.065 59.150 ;
        RECT 143.820 58.890 144.080 59.150 ;
        RECT 144.140 58.890 144.400 59.150 ;
        RECT 144.460 58.890 144.720 59.150 ;
        RECT 144.780 58.890 145.040 59.150 ;
        RECT 145.100 58.890 145.360 59.150 ;
        RECT 96.680 58.380 96.940 58.640 ;
        RECT 97.600 57.360 97.860 57.620 ;
        RECT 99.900 58.380 100.160 58.640 ;
        RECT 100.820 58.380 101.080 58.640 ;
        RECT 107.260 58.380 107.520 58.640 ;
        RECT 110.940 58.380 111.200 58.640 ;
        RECT 150.040 58.380 150.300 58.640 ;
        RECT 98.980 57.360 99.240 57.620 ;
        RECT 131.180 57.700 131.440 57.960 ;
        RECT 142.680 57.700 142.940 57.960 ;
        RECT 100.360 57.360 100.620 57.620 ;
        RECT 102.200 57.360 102.460 57.620 ;
        RECT 120.600 57.360 120.860 57.620 ;
        RECT 123.820 57.360 124.080 57.620 ;
        RECT 126.120 57.360 126.380 57.620 ;
        RECT 127.960 57.360 128.220 57.620 ;
        RECT 135.320 57.360 135.580 57.620 ;
        RECT 141.300 57.360 141.560 57.620 ;
        RECT 97.140 57.020 97.400 57.280 ;
        RECT 130.260 57.020 130.520 57.280 ;
        RECT 136.240 57.020 136.500 57.280 ;
        RECT 147.740 57.020 148.000 57.280 ;
        RECT 96.680 56.680 96.940 56.940 ;
        RECT 118.300 56.680 118.560 56.940 ;
        RECT 125.660 56.680 125.920 56.940 ;
        RECT 127.500 56.680 127.760 56.940 ;
        RECT 133.480 56.680 133.740 56.940 ;
        RECT 101.235 56.170 101.495 56.430 ;
        RECT 101.555 56.170 101.815 56.430 ;
        RECT 101.875 56.170 102.135 56.430 ;
        RECT 102.195 56.170 102.455 56.430 ;
        RECT 102.515 56.170 102.775 56.430 ;
        RECT 116.530 56.170 116.790 56.430 ;
        RECT 116.850 56.170 117.110 56.430 ;
        RECT 117.170 56.170 117.430 56.430 ;
        RECT 117.490 56.170 117.750 56.430 ;
        RECT 117.810 56.170 118.070 56.430 ;
        RECT 131.825 56.170 132.085 56.430 ;
        RECT 132.145 56.170 132.405 56.430 ;
        RECT 132.465 56.170 132.725 56.430 ;
        RECT 132.785 56.170 133.045 56.430 ;
        RECT 133.105 56.170 133.365 56.430 ;
        RECT 147.120 56.170 147.380 56.430 ;
        RECT 147.440 56.170 147.700 56.430 ;
        RECT 147.760 56.170 148.020 56.430 ;
        RECT 148.080 56.170 148.340 56.430 ;
        RECT 148.400 56.170 148.660 56.430 ;
        RECT 97.600 55.660 97.860 55.920 ;
        RECT 98.980 54.980 99.240 55.240 ;
        RECT 100.360 54.980 100.620 55.240 ;
        RECT 103.120 54.980 103.380 55.240 ;
        RECT 115.080 54.980 115.340 55.240 ;
        RECT 127.500 55.660 127.760 55.920 ;
        RECT 118.300 54.980 118.560 55.240 ;
        RECT 125.660 55.320 125.920 55.580 ;
        RECT 130.720 54.980 130.980 55.240 ;
        RECT 133.480 55.320 133.740 55.580 ;
        RECT 141.300 55.320 141.560 55.580 ;
        RECT 145.900 54.980 146.160 55.240 ;
        RECT 142.680 54.640 142.940 54.900 ;
        RECT 110.480 54.300 110.740 54.560 ;
        RECT 108.640 53.960 108.900 54.220 ;
        RECT 115.540 53.960 115.800 54.220 ;
        RECT 118.300 53.960 118.560 54.220 ;
        RECT 120.140 53.960 120.400 54.220 ;
        RECT 121.980 53.960 122.240 54.220 ;
        RECT 136.240 53.960 136.500 54.220 ;
        RECT 147.740 53.960 148.000 54.220 ;
        RECT 97.935 53.450 98.195 53.710 ;
        RECT 98.255 53.450 98.515 53.710 ;
        RECT 98.575 53.450 98.835 53.710 ;
        RECT 98.895 53.450 99.155 53.710 ;
        RECT 99.215 53.450 99.475 53.710 ;
        RECT 113.230 53.450 113.490 53.710 ;
        RECT 113.550 53.450 113.810 53.710 ;
        RECT 113.870 53.450 114.130 53.710 ;
        RECT 114.190 53.450 114.450 53.710 ;
        RECT 114.510 53.450 114.770 53.710 ;
        RECT 128.525 53.450 128.785 53.710 ;
        RECT 128.845 53.450 129.105 53.710 ;
        RECT 129.165 53.450 129.425 53.710 ;
        RECT 129.485 53.450 129.745 53.710 ;
        RECT 129.805 53.450 130.065 53.710 ;
        RECT 143.820 53.450 144.080 53.710 ;
        RECT 144.140 53.450 144.400 53.710 ;
        RECT 144.460 53.450 144.720 53.710 ;
        RECT 144.780 53.450 145.040 53.710 ;
        RECT 145.100 53.450 145.360 53.710 ;
        RECT 96.680 52.940 96.940 53.200 ;
        RECT 115.540 52.940 115.800 53.200 ;
        RECT 118.300 52.940 118.560 53.200 ;
        RECT 127.960 52.940 128.220 53.200 ;
        RECT 133.480 52.940 133.740 53.200 ;
        RECT 140.380 52.940 140.640 53.200 ;
        RECT 106.340 52.260 106.600 52.520 ;
        RECT 92.540 51.920 92.800 52.180 ;
        RECT 100.820 51.920 101.080 52.180 ;
        RECT 103.120 51.920 103.380 52.180 ;
        RECT 110.020 51.920 110.280 52.180 ;
        RECT 110.940 52.260 111.200 52.520 ;
        RECT 112.780 52.260 113.040 52.520 ;
        RECT 135.320 52.260 135.580 52.520 ;
        RECT 137.620 52.260 137.880 52.520 ;
        RECT 111.400 51.920 111.660 52.180 ;
        RECT 120.140 51.920 120.400 52.180 ;
        RECT 121.980 51.920 122.240 52.180 ;
        RECT 104.040 51.580 104.300 51.840 ;
        RECT 106.800 51.580 107.060 51.840 ;
        RECT 107.720 51.580 107.980 51.840 ;
        RECT 112.320 51.580 112.580 51.840 ;
        RECT 115.080 51.580 115.340 51.840 ;
        RECT 121.520 51.580 121.780 51.840 ;
        RECT 130.260 51.920 130.520 52.180 ;
        RECT 130.720 51.920 130.980 52.180 ;
        RECT 131.180 51.920 131.440 52.180 ;
        RECT 100.360 51.240 100.620 51.500 ;
        RECT 108.180 51.240 108.440 51.500 ;
        RECT 109.100 51.240 109.360 51.500 ;
        RECT 122.440 51.240 122.700 51.500 ;
        RECT 127.500 51.240 127.760 51.500 ;
        RECT 134.400 51.920 134.660 52.180 ;
        RECT 134.860 51.920 135.120 52.180 ;
        RECT 134.400 51.240 134.660 51.500 ;
        RECT 136.240 51.580 136.500 51.840 ;
        RECT 138.540 51.240 138.800 51.500 ;
        RECT 141.300 51.920 141.560 52.180 ;
        RECT 147.740 51.580 148.000 51.840 ;
        RECT 101.235 50.730 101.495 50.990 ;
        RECT 101.555 50.730 101.815 50.990 ;
        RECT 101.875 50.730 102.135 50.990 ;
        RECT 102.195 50.730 102.455 50.990 ;
        RECT 102.515 50.730 102.775 50.990 ;
        RECT 116.530 50.730 116.790 50.990 ;
        RECT 116.850 50.730 117.110 50.990 ;
        RECT 117.170 50.730 117.430 50.990 ;
        RECT 117.490 50.730 117.750 50.990 ;
        RECT 117.810 50.730 118.070 50.990 ;
        RECT 131.825 50.730 132.085 50.990 ;
        RECT 132.145 50.730 132.405 50.990 ;
        RECT 132.465 50.730 132.725 50.990 ;
        RECT 132.785 50.730 133.045 50.990 ;
        RECT 133.105 50.730 133.365 50.990 ;
        RECT 147.120 50.730 147.380 50.990 ;
        RECT 147.440 50.730 147.700 50.990 ;
        RECT 147.760 50.730 148.020 50.990 ;
        RECT 148.080 50.730 148.340 50.990 ;
        RECT 148.400 50.730 148.660 50.990 ;
        RECT 107.720 50.220 107.980 50.480 ;
        RECT 109.100 50.220 109.360 50.480 ;
        RECT 110.480 50.220 110.740 50.480 ;
        RECT 121.520 50.220 121.780 50.480 ;
        RECT 127.500 50.220 127.760 50.480 ;
        RECT 128.880 50.220 129.140 50.480 ;
        RECT 133.940 50.220 134.200 50.480 ;
        RECT 134.400 50.220 134.660 50.480 ;
        RECT 92.540 49.880 92.800 50.140 ;
        RECT 97.140 49.200 97.400 49.460 ;
        RECT 101.280 49.540 101.540 49.800 ;
        RECT 100.820 49.200 101.080 49.460 ;
        RECT 106.800 49.880 107.060 50.140 ;
        RECT 104.040 49.200 104.300 49.460 ;
        RECT 105.880 49.200 106.140 49.460 ;
        RECT 115.080 49.880 115.340 50.140 ;
        RECT 121.980 49.880 122.240 50.140 ;
        RECT 131.180 49.880 131.440 50.140 ;
        RECT 106.800 49.200 107.060 49.460 ;
        RECT 111.860 49.200 112.120 49.460 ;
        RECT 133.480 49.540 133.740 49.800 ;
        RECT 134.860 49.880 135.120 50.140 ;
        RECT 135.780 50.220 136.040 50.480 ;
        RECT 138.540 50.220 138.800 50.480 ;
        RECT 128.880 49.200 129.140 49.460 ;
        RECT 134.400 49.200 134.660 49.460 ;
        RECT 137.620 49.880 137.880 50.140 ;
        RECT 145.440 49.540 145.700 49.800 ;
        RECT 150.500 49.200 150.760 49.460 ;
        RECT 96.220 48.520 96.480 48.780 ;
        RECT 99.900 48.520 100.160 48.780 ;
        RECT 105.420 48.520 105.680 48.780 ;
        RECT 110.940 48.520 111.200 48.780 ;
        RECT 97.935 48.010 98.195 48.270 ;
        RECT 98.255 48.010 98.515 48.270 ;
        RECT 98.575 48.010 98.835 48.270 ;
        RECT 98.895 48.010 99.155 48.270 ;
        RECT 99.215 48.010 99.475 48.270 ;
        RECT 113.230 48.010 113.490 48.270 ;
        RECT 113.550 48.010 113.810 48.270 ;
        RECT 113.870 48.010 114.130 48.270 ;
        RECT 114.190 48.010 114.450 48.270 ;
        RECT 114.510 48.010 114.770 48.270 ;
        RECT 128.525 48.010 128.785 48.270 ;
        RECT 128.845 48.010 129.105 48.270 ;
        RECT 129.165 48.010 129.425 48.270 ;
        RECT 129.485 48.010 129.745 48.270 ;
        RECT 129.805 48.010 130.065 48.270 ;
        RECT 143.820 48.010 144.080 48.270 ;
        RECT 144.140 48.010 144.400 48.270 ;
        RECT 144.460 48.010 144.720 48.270 ;
        RECT 144.780 48.010 145.040 48.270 ;
        RECT 145.100 48.010 145.360 48.270 ;
        RECT 92.540 47.500 92.800 47.760 ;
        RECT 107.260 47.500 107.520 47.760 ;
        RECT 107.720 47.500 107.980 47.760 ;
        RECT 108.180 47.500 108.440 47.760 ;
        RECT 110.020 47.500 110.280 47.760 ;
        RECT 110.940 47.500 111.200 47.760 ;
        RECT 111.400 47.500 111.660 47.760 ;
        RECT 120.140 47.500 120.400 47.760 ;
        RECT 96.220 46.820 96.480 47.080 ;
        RECT 99.900 46.480 100.160 46.740 ;
        RECT 105.420 45.800 105.680 46.060 ;
        RECT 129.340 47.160 129.600 47.420 ;
        RECT 130.720 46.820 130.980 47.080 ;
        RECT 120.600 45.800 120.860 46.060 ;
        RECT 126.580 46.140 126.840 46.400 ;
        RECT 101.235 45.290 101.495 45.550 ;
        RECT 101.555 45.290 101.815 45.550 ;
        RECT 101.875 45.290 102.135 45.550 ;
        RECT 102.195 45.290 102.455 45.550 ;
        RECT 102.515 45.290 102.775 45.550 ;
        RECT 116.530 45.290 116.790 45.550 ;
        RECT 116.850 45.290 117.110 45.550 ;
        RECT 117.170 45.290 117.430 45.550 ;
        RECT 117.490 45.290 117.750 45.550 ;
        RECT 117.810 45.290 118.070 45.550 ;
        RECT 131.825 45.290 132.085 45.550 ;
        RECT 132.145 45.290 132.405 45.550 ;
        RECT 132.465 45.290 132.725 45.550 ;
        RECT 132.785 45.290 133.045 45.550 ;
        RECT 133.105 45.290 133.365 45.550 ;
        RECT 147.120 45.290 147.380 45.550 ;
        RECT 147.440 45.290 147.700 45.550 ;
        RECT 147.760 45.290 148.020 45.550 ;
        RECT 148.080 45.290 148.340 45.550 ;
        RECT 148.400 45.290 148.660 45.550 ;
        RECT 100.820 44.780 101.080 45.040 ;
        RECT 110.480 44.780 110.740 45.040 ;
        RECT 111.860 44.780 112.120 45.040 ;
        RECT 115.080 44.780 115.340 45.040 ;
        RECT 129.340 44.780 129.600 45.040 ;
        RECT 131.180 44.780 131.440 45.040 ;
        RECT 134.400 44.780 134.660 45.040 ;
        RECT 134.860 44.780 135.120 45.040 ;
        RECT 97.140 44.440 97.400 44.700 ;
        RECT 105.880 44.440 106.140 44.700 ;
        RECT 113.240 44.440 113.500 44.700 ;
        RECT 127.040 44.440 127.300 44.700 ;
        RECT 104.040 44.100 104.300 44.360 ;
        RECT 105.420 44.100 105.680 44.360 ;
        RECT 120.140 44.100 120.400 44.360 ;
        RECT 127.040 43.760 127.300 44.020 ;
        RECT 127.960 44.100 128.220 44.360 ;
        RECT 131.640 44.100 131.900 44.360 ;
        RECT 139.000 44.440 139.260 44.700 ;
        RECT 140.840 44.440 141.100 44.700 ;
        RECT 134.860 43.760 135.120 44.020 ;
        RECT 142.680 43.760 142.940 44.020 ;
        RECT 96.220 43.080 96.480 43.340 ;
        RECT 107.260 43.080 107.520 43.340 ;
        RECT 126.580 43.080 126.840 43.340 ;
        RECT 134.400 43.080 134.660 43.340 ;
        RECT 141.760 43.080 142.020 43.340 ;
        RECT 143.140 43.080 143.400 43.340 ;
        RECT 146.360 43.080 146.620 43.340 ;
        RECT 97.935 42.570 98.195 42.830 ;
        RECT 98.255 42.570 98.515 42.830 ;
        RECT 98.575 42.570 98.835 42.830 ;
        RECT 98.895 42.570 99.155 42.830 ;
        RECT 99.215 42.570 99.475 42.830 ;
        RECT 113.230 42.570 113.490 42.830 ;
        RECT 113.550 42.570 113.810 42.830 ;
        RECT 113.870 42.570 114.130 42.830 ;
        RECT 114.190 42.570 114.450 42.830 ;
        RECT 114.510 42.570 114.770 42.830 ;
        RECT 128.525 42.570 128.785 42.830 ;
        RECT 128.845 42.570 129.105 42.830 ;
        RECT 129.165 42.570 129.425 42.830 ;
        RECT 129.485 42.570 129.745 42.830 ;
        RECT 129.805 42.570 130.065 42.830 ;
        RECT 143.820 42.570 144.080 42.830 ;
        RECT 144.140 42.570 144.400 42.830 ;
        RECT 144.460 42.570 144.720 42.830 ;
        RECT 144.780 42.570 145.040 42.830 ;
        RECT 145.100 42.570 145.360 42.830 ;
        RECT 131.640 42.060 131.900 42.320 ;
        RECT 142.680 42.060 142.940 42.320 ;
        RECT 149.580 42.060 149.840 42.320 ;
        RECT 109.560 41.380 109.820 41.640 ;
        RECT 143.140 41.380 143.400 41.640 ;
        RECT 90.240 41.040 90.500 41.300 ;
        RECT 96.220 40.360 96.480 40.620 ;
        RECT 139.000 41.040 139.260 41.300 ;
        RECT 140.380 40.700 140.640 40.960 ;
        RECT 141.300 41.040 141.560 41.300 ;
        RECT 146.360 40.700 146.620 40.960 ;
        RECT 140.840 40.360 141.100 40.620 ;
        RECT 142.220 40.360 142.480 40.620 ;
        RECT 101.235 39.850 101.495 40.110 ;
        RECT 101.555 39.850 101.815 40.110 ;
        RECT 101.875 39.850 102.135 40.110 ;
        RECT 102.195 39.850 102.455 40.110 ;
        RECT 102.515 39.850 102.775 40.110 ;
        RECT 116.530 39.850 116.790 40.110 ;
        RECT 116.850 39.850 117.110 40.110 ;
        RECT 117.170 39.850 117.430 40.110 ;
        RECT 117.490 39.850 117.750 40.110 ;
        RECT 117.810 39.850 118.070 40.110 ;
        RECT 131.825 39.850 132.085 40.110 ;
        RECT 132.145 39.850 132.405 40.110 ;
        RECT 132.465 39.850 132.725 40.110 ;
        RECT 132.785 39.850 133.045 40.110 ;
        RECT 133.105 39.850 133.365 40.110 ;
        RECT 147.120 39.850 147.380 40.110 ;
        RECT 147.440 39.850 147.700 40.110 ;
        RECT 147.760 39.850 148.020 40.110 ;
        RECT 148.080 39.850 148.340 40.110 ;
        RECT 148.400 39.850 148.660 40.110 ;
        RECT 1.280 35.295 2.220 36.155 ;
        RECT 102.200 39.340 102.460 39.600 ;
        RECT 106.340 39.340 106.600 39.600 ;
        RECT 95.760 38.320 96.020 38.580 ;
        RECT 96.680 38.320 96.940 38.580 ;
        RECT 98.980 38.320 99.240 38.580 ;
        RECT 107.260 38.660 107.520 38.920 ;
        RECT 104.040 38.320 104.300 38.580 ;
        RECT 115.540 39.000 115.800 39.260 ;
        RECT 109.560 38.660 109.820 38.920 ;
        RECT 110.020 38.660 110.280 38.920 ;
        RECT 121.520 39.340 121.780 39.600 ;
        RECT 121.980 39.340 122.240 39.600 ;
        RECT 122.440 38.660 122.700 38.920 ;
        RECT 123.360 38.660 123.620 38.920 ;
        RECT 124.280 38.660 124.540 38.920 ;
        RECT 100.820 37.980 101.080 38.240 ;
        RECT 103.580 37.980 103.840 38.240 ;
        RECT 105.420 37.980 105.680 38.240 ;
        RECT 112.320 38.320 112.580 38.580 ;
        RECT 115.080 38.320 115.340 38.580 ;
        RECT 116.000 38.320 116.260 38.580 ;
        RECT 117.840 38.320 118.100 38.580 ;
        RECT 119.680 38.320 119.940 38.580 ;
        RECT 125.660 38.660 125.920 38.920 ;
        RECT 126.120 38.660 126.380 38.920 ;
        RECT 127.500 38.660 127.760 38.920 ;
        RECT 111.860 37.980 112.120 38.240 ;
        RECT 112.780 37.980 113.040 38.240 ;
        RECT 121.060 37.980 121.320 38.240 ;
        RECT 121.520 37.980 121.780 38.240 ;
        RECT 139.920 39.340 140.180 39.600 ;
        RECT 140.380 39.340 140.640 39.600 ;
        RECT 142.220 39.340 142.480 39.600 ;
        RECT 140.840 39.000 141.100 39.260 ;
        RECT 134.400 38.660 134.660 38.920 ;
        RECT 134.860 38.660 135.120 38.920 ;
        RECT 139.920 38.660 140.180 38.920 ;
        RECT 150.040 38.660 150.300 38.920 ;
        RECT 139.000 38.320 139.260 38.580 ;
        RECT 99.900 37.640 100.160 37.900 ;
        RECT 104.960 37.640 105.220 37.900 ;
        RECT 110.940 37.640 111.200 37.900 ;
        RECT 111.400 37.640 111.660 37.900 ;
        RECT 118.760 37.640 119.020 37.900 ;
        RECT 120.140 37.640 120.400 37.900 ;
        RECT 123.360 37.640 123.620 37.900 ;
        RECT 131.180 37.980 131.440 38.240 ;
        RECT 131.640 37.980 131.900 38.240 ;
        RECT 127.500 37.640 127.760 37.900 ;
        RECT 127.960 37.640 128.220 37.900 ;
        RECT 130.260 37.640 130.520 37.900 ;
        RECT 130.720 37.640 130.980 37.900 ;
        RECT 137.620 37.980 137.880 38.240 ;
        RECT 141.760 38.320 142.020 38.580 ;
        RECT 139.460 37.640 139.720 37.900 ;
        RECT 145.900 37.640 146.160 37.900 ;
        RECT 97.935 37.130 98.195 37.390 ;
        RECT 98.255 37.130 98.515 37.390 ;
        RECT 98.575 37.130 98.835 37.390 ;
        RECT 98.895 37.130 99.155 37.390 ;
        RECT 99.215 37.130 99.475 37.390 ;
        RECT 113.230 37.130 113.490 37.390 ;
        RECT 113.550 37.130 113.810 37.390 ;
        RECT 113.870 37.130 114.130 37.390 ;
        RECT 114.190 37.130 114.450 37.390 ;
        RECT 114.510 37.130 114.770 37.390 ;
        RECT 128.525 37.130 128.785 37.390 ;
        RECT 128.845 37.130 129.105 37.390 ;
        RECT 129.165 37.130 129.425 37.390 ;
        RECT 129.485 37.130 129.745 37.390 ;
        RECT 129.805 37.130 130.065 37.390 ;
        RECT 143.820 37.130 144.080 37.390 ;
        RECT 144.140 37.130 144.400 37.390 ;
        RECT 144.460 37.130 144.720 37.390 ;
        RECT 144.780 37.130 145.040 37.390 ;
        RECT 145.100 37.130 145.360 37.390 ;
        RECT 93.460 35.600 93.720 35.860 ;
        RECT 96.680 36.280 96.940 36.540 ;
        RECT 95.760 35.940 96.020 36.200 ;
        RECT 99.900 36.620 100.160 36.880 ;
        RECT 100.360 35.940 100.620 36.200 ;
        RECT 100.820 35.600 101.080 35.860 ;
        RECT 102.200 36.280 102.460 36.540 ;
        RECT 103.580 35.600 103.840 35.860 ;
        RECT 105.880 35.940 106.140 36.200 ;
        RECT 109.560 36.620 109.820 36.880 ;
        RECT 110.940 36.620 111.200 36.880 ;
        RECT 119.680 36.620 119.940 36.880 ;
        RECT 116.000 36.280 116.260 36.540 ;
        RECT 112.780 35.940 113.040 36.200 ;
        RECT 115.540 35.940 115.800 36.200 ;
        RECT 120.140 36.280 120.400 36.540 ;
        RECT 121.060 36.620 121.320 36.880 ;
        RECT 125.660 36.620 125.920 36.880 ;
        RECT 107.260 35.600 107.520 35.860 ;
        RECT 109.560 35.600 109.820 35.860 ;
        RECT 95.760 34.920 96.020 35.180 ;
        RECT 99.900 34.920 100.160 35.180 ;
        RECT 110.940 35.600 111.200 35.860 ;
        RECT 111.860 35.600 112.120 35.860 ;
        RECT 116.000 35.600 116.260 35.860 ;
        RECT 114.620 34.920 114.880 35.180 ;
        RECT 119.220 35.600 119.480 35.860 ;
        RECT 121.060 35.940 121.320 36.200 ;
        RECT 121.980 35.940 122.240 36.200 ;
        RECT 120.140 35.260 120.400 35.520 ;
        RECT 121.520 35.600 121.780 35.860 ;
        RECT 124.280 35.940 124.540 36.200 ;
        RECT 127.960 35.940 128.220 36.200 ;
        RECT 129.800 35.940 130.060 36.200 ;
        RECT 131.640 36.620 131.900 36.880 ;
        RECT 139.000 36.620 139.260 36.880 ;
        RECT 139.920 36.620 140.180 36.880 ;
        RECT 150.040 36.620 150.300 36.880 ;
        RECT 126.580 35.600 126.840 35.860 ;
        RECT 127.500 35.600 127.760 35.860 ;
        RECT 128.420 35.600 128.680 35.860 ;
        RECT 128.880 35.600 129.140 35.860 ;
        RECT 130.720 35.600 130.980 35.860 ;
        RECT 132.560 36.280 132.820 36.540 ;
        RECT 133.480 36.280 133.740 36.540 ;
        RECT 134.400 36.280 134.660 36.540 ;
        RECT 132.100 35.600 132.360 35.860 ;
        RECT 133.480 35.600 133.740 35.860 ;
        RECT 133.940 35.600 134.200 35.860 ;
        RECT 134.400 35.600 134.660 35.860 ;
        RECT 141.300 35.940 141.560 36.200 ;
        RECT 122.900 34.920 123.160 35.180 ;
        RECT 126.580 34.920 126.840 35.180 ;
        RECT 127.040 34.920 127.300 35.180 ;
        RECT 130.260 35.260 130.520 35.520 ;
        RECT 130.720 34.920 130.980 35.180 ;
        RECT 132.100 34.920 132.360 35.180 ;
        RECT 132.560 34.920 132.820 35.180 ;
        RECT 139.920 35.600 140.180 35.860 ;
        RECT 140.380 35.600 140.640 35.860 ;
        RECT 140.840 34.920 141.100 35.180 ;
        RECT 149.120 35.260 149.380 35.520 ;
        RECT 146.360 34.920 146.620 35.180 ;
        RECT 101.235 34.410 101.495 34.670 ;
        RECT 101.555 34.410 101.815 34.670 ;
        RECT 101.875 34.410 102.135 34.670 ;
        RECT 102.195 34.410 102.455 34.670 ;
        RECT 102.515 34.410 102.775 34.670 ;
        RECT 116.530 34.410 116.790 34.670 ;
        RECT 116.850 34.410 117.110 34.670 ;
        RECT 117.170 34.410 117.430 34.670 ;
        RECT 117.490 34.410 117.750 34.670 ;
        RECT 117.810 34.410 118.070 34.670 ;
        RECT 131.825 34.410 132.085 34.670 ;
        RECT 132.145 34.410 132.405 34.670 ;
        RECT 132.465 34.410 132.725 34.670 ;
        RECT 132.785 34.410 133.045 34.670 ;
        RECT 133.105 34.410 133.365 34.670 ;
        RECT 147.120 34.410 147.380 34.670 ;
        RECT 147.440 34.410 147.700 34.670 ;
        RECT 147.760 34.410 148.020 34.670 ;
        RECT 148.080 34.410 148.340 34.670 ;
        RECT 148.400 34.410 148.660 34.670 ;
        RECT 8.050 28.940 8.415 29.470 ;
        RECT 99.900 33.900 100.160 34.160 ;
        RECT 100.820 33.900 101.080 34.160 ;
        RECT 102.200 33.900 102.460 34.160 ;
        RECT 104.960 33.900 105.220 34.160 ;
        RECT 105.880 33.900 106.140 34.160 ;
        RECT 106.340 33.900 106.600 34.160 ;
        RECT 99.900 33.220 100.160 33.480 ;
        RECT 102.660 33.220 102.920 33.480 ;
        RECT 104.040 33.220 104.300 33.480 ;
        RECT 105.880 33.220 106.140 33.480 ;
        RECT 110.020 33.900 110.280 34.160 ;
        RECT 111.400 33.900 111.660 34.160 ;
        RECT 115.080 33.900 115.340 34.160 ;
        RECT 118.760 33.900 119.020 34.160 ;
        RECT 120.140 33.900 120.400 34.160 ;
        RECT 124.280 33.900 124.540 34.160 ;
        RECT 126.120 33.900 126.380 34.160 ;
        RECT 126.580 33.900 126.840 34.160 ;
        RECT 116.000 33.560 116.260 33.820 ;
        RECT 128.420 33.900 128.680 34.160 ;
        RECT 131.180 33.900 131.440 34.160 ;
        RECT 107.720 32.880 107.980 33.140 ;
        RECT 111.400 33.220 111.660 33.480 ;
        RECT 112.320 33.220 112.580 33.480 ;
        RECT 112.780 33.220 113.040 33.480 ;
        RECT 114.620 33.220 114.880 33.480 ;
        RECT 115.540 33.220 115.800 33.480 ;
        RECT 117.840 33.220 118.100 33.480 ;
        RECT 122.900 33.220 123.160 33.480 ;
        RECT 127.040 33.220 127.300 33.480 ;
        RECT 127.960 33.220 128.220 33.480 ;
        RECT 130.260 33.220 130.520 33.480 ;
        RECT 132.100 33.560 132.360 33.820 ;
        RECT 133.940 33.900 134.200 34.160 ;
        RECT 146.360 33.900 146.620 34.160 ;
        RECT 149.120 33.900 149.380 34.160 ;
        RECT 149.580 33.900 149.840 34.160 ;
        RECT 137.620 33.560 137.880 33.820 ;
        RECT 134.400 33.220 134.660 33.480 ;
        RECT 145.900 33.220 146.160 33.480 ;
        RECT 152.800 33.220 153.060 33.480 ;
        RECT 102.200 32.200 102.460 32.460 ;
        RECT 105.420 32.540 105.680 32.800 ;
        RECT 105.880 32.540 106.140 32.800 ;
        RECT 109.560 32.540 109.820 32.800 ;
        RECT 137.620 32.880 137.880 33.140 ;
        RECT 139.920 32.880 140.180 33.140 ;
        RECT 127.500 32.540 127.760 32.800 ;
        RECT 140.840 32.540 141.100 32.800 ;
        RECT 110.940 32.200 111.200 32.460 ;
        RECT 111.400 32.200 111.660 32.460 ;
        RECT 97.935 31.690 98.195 31.950 ;
        RECT 98.255 31.690 98.515 31.950 ;
        RECT 98.575 31.690 98.835 31.950 ;
        RECT 98.895 31.690 99.155 31.950 ;
        RECT 99.215 31.690 99.475 31.950 ;
        RECT 113.230 31.690 113.490 31.950 ;
        RECT 113.550 31.690 113.810 31.950 ;
        RECT 113.870 31.690 114.130 31.950 ;
        RECT 114.190 31.690 114.450 31.950 ;
        RECT 114.510 31.690 114.770 31.950 ;
        RECT 128.525 31.690 128.785 31.950 ;
        RECT 128.845 31.690 129.105 31.950 ;
        RECT 129.165 31.690 129.425 31.950 ;
        RECT 129.485 31.690 129.745 31.950 ;
        RECT 129.805 31.690 130.065 31.950 ;
        RECT 143.820 31.690 144.080 31.950 ;
        RECT 144.140 31.690 144.400 31.950 ;
        RECT 144.460 31.690 144.720 31.950 ;
        RECT 144.780 31.690 145.040 31.950 ;
        RECT 145.100 31.690 145.360 31.950 ;
        RECT 93.460 31.180 93.720 31.440 ;
        RECT 99.900 31.180 100.160 31.440 ;
        RECT 107.720 31.180 107.980 31.440 ;
        RECT 111.400 31.180 111.660 31.440 ;
        RECT 115.540 31.180 115.800 31.440 ;
        RECT 117.840 31.180 118.100 31.440 ;
        RECT 130.260 31.180 130.520 31.440 ;
        RECT 137.620 31.180 137.880 31.440 ;
        RECT 150.960 31.180 151.220 31.440 ;
        RECT 90.240 30.160 90.500 30.420 ;
        RECT 98.520 30.160 98.780 30.420 ;
        RECT 106.340 30.160 106.600 30.420 ;
        RECT 114.160 30.160 114.420 30.420 ;
        RECT 116.000 30.160 116.260 30.420 ;
        RECT 140.840 30.500 141.100 30.760 ;
        RECT 121.520 30.160 121.780 30.420 ;
        RECT 129.340 30.160 129.600 30.420 ;
        RECT 137.160 30.160 137.420 30.420 ;
        RECT 144.980 29.820 145.240 30.080 ;
        RECT 151.880 29.820 152.140 30.080 ;
        RECT 101.235 28.970 101.495 29.230 ;
        RECT 101.555 28.970 101.815 29.230 ;
        RECT 101.875 28.970 102.135 29.230 ;
        RECT 102.195 28.970 102.455 29.230 ;
        RECT 102.515 28.970 102.775 29.230 ;
        RECT 116.530 28.970 116.790 29.230 ;
        RECT 116.850 28.970 117.110 29.230 ;
        RECT 117.170 28.970 117.430 29.230 ;
        RECT 117.490 28.970 117.750 29.230 ;
        RECT 117.810 28.970 118.070 29.230 ;
        RECT 131.825 28.970 132.085 29.230 ;
        RECT 132.145 28.970 132.405 29.230 ;
        RECT 132.465 28.970 132.725 29.230 ;
        RECT 132.785 28.970 133.045 29.230 ;
        RECT 133.105 28.970 133.365 29.230 ;
        RECT 147.120 28.970 147.380 29.230 ;
        RECT 147.440 28.970 147.700 29.230 ;
        RECT 147.760 28.970 148.020 29.230 ;
        RECT 148.080 28.970 148.340 29.230 ;
        RECT 148.400 28.970 148.660 29.230 ;
        RECT 1.280 23.810 2.220 24.670 ;
        RECT 59.095 20.600 59.375 20.880 ;
        RECT 8.560 16.620 9.610 17.985 ;
        RECT 53.335 8.005 53.805 8.460 ;
        RECT 83.210 7.760 83.645 8.180 ;
      LAYER met2 ;
        RECT 84.935 222.850 85.235 222.915 ;
        RECT 84.925 222.590 85.245 222.850 ;
        RECT 84.935 222.525 85.235 222.590 ;
        RECT 88.605 222.530 88.905 222.920 ;
        RECT 4.955 211.625 5.675 211.770 ;
        RECT 88.615 211.625 88.895 222.530 ;
        RECT 157.210 221.425 157.855 221.455 ;
        RECT 147.305 220.825 157.855 221.425 ;
        RECT 157.210 220.800 157.855 220.825 ;
        RECT 143.605 219.560 144.325 219.620 ;
        RECT 155.965 219.560 156.615 219.590 ;
        RECT 143.605 218.960 156.615 219.560 ;
        RECT 143.605 218.905 144.325 218.960 ;
        RECT 155.965 218.935 156.615 218.960 ;
        RECT 139.920 217.380 140.640 217.440 ;
        RECT 153.605 217.380 154.255 217.405 ;
        RECT 139.920 216.780 154.255 217.380 ;
        RECT 139.920 216.725 140.640 216.780 ;
        RECT 153.605 216.750 154.255 216.780 ;
        RECT 136.265 215.715 136.985 215.770 ;
        RECT 153.840 215.715 154.490 215.745 ;
        RECT 136.265 215.115 154.490 215.715 ;
        RECT 136.265 215.055 136.985 215.115 ;
        RECT 153.840 215.090 154.490 215.115 ;
        RECT 4.955 211.345 110.720 211.625 ;
        RECT 4.955 211.330 5.675 211.345 ;
        RECT 3.475 207.765 4.045 207.825 ;
        RECT 80.540 207.765 80.820 207.800 ;
        RECT 3.475 207.485 80.820 207.765 ;
        RECT 3.475 207.405 4.045 207.485 ;
        RECT 80.540 203.800 80.820 207.485 ;
        RECT 110.440 203.800 110.720 211.345 ;
        RECT 80.610 200.510 80.750 203.800 ;
        RECT 84.950 200.510 85.210 200.595 ;
        RECT 80.600 200.355 85.210 200.510 ;
        RECT 1.005 193.685 2.505 195.185 ;
        RECT 76.515 194.245 78.055 194.615 ;
        RECT 80.610 194.080 80.750 200.355 ;
        RECT 84.950 200.275 85.210 200.355 ;
        RECT 88.590 194.245 90.130 194.615 ;
        RECT 100.665 194.245 102.205 194.615 ;
        RECT 110.510 194.080 110.650 203.800 ;
        RECT 112.740 194.245 114.280 194.615 ;
        RECT 80.550 193.760 80.810 194.080 ;
        RECT 110.450 193.760 110.710 194.080 ;
        RECT 86.990 192.740 87.250 193.060 ;
        RECT 81.470 192.400 81.730 192.720 ;
        RECT 79.815 191.525 81.355 191.895 ;
        RECT 81.530 191.360 81.670 192.400 ;
        RECT 82.390 192.060 82.650 192.380 ;
        RECT 81.470 191.040 81.730 191.360 ;
        RECT 70.430 190.360 70.690 190.680 ;
        RECT 81.010 190.360 81.270 190.680 ;
        RECT 70.490 189.515 70.630 190.360 ;
        RECT 70.420 189.145 70.700 189.515 ;
        RECT 73.650 189.340 73.910 189.660 ;
        RECT 73.710 188.640 73.850 189.340 ;
        RECT 76.515 188.805 78.055 189.175 ;
        RECT 73.650 188.320 73.910 188.640 ;
        RECT 81.070 186.850 81.210 190.360 ;
        RECT 82.450 188.640 82.590 192.060 ;
        RECT 82.850 190.360 83.110 190.680 ;
        RECT 82.910 188.640 83.050 190.360 ;
        RECT 83.770 189.680 84.030 190.000 ;
        RECT 82.390 188.320 82.650 188.640 ;
        RECT 82.850 188.320 83.110 188.640 ;
        RECT 83.830 187.620 83.970 189.680 ;
        RECT 87.050 189.660 87.190 192.740 ;
        RECT 100.330 192.400 100.590 192.720 ;
        RECT 102.630 192.400 102.890 192.720 ;
        RECT 111.370 192.400 111.630 192.720 ;
        RECT 91.890 191.525 93.430 191.895 ;
        RECT 100.390 190.680 100.530 192.400 ;
        RECT 100.330 190.360 100.590 190.680 ;
        RECT 87.910 190.020 88.170 190.340 ;
        RECT 94.810 190.020 95.070 190.340 ;
        RECT 84.230 189.340 84.490 189.660 ;
        RECT 86.990 189.340 87.250 189.660 ;
        RECT 83.770 187.300 84.030 187.620 ;
        RECT 81.070 186.710 82.130 186.850 ;
        RECT 79.815 186.085 81.355 186.455 ;
        RECT 79.170 185.600 79.430 185.920 ;
        RECT 76.515 183.365 78.055 183.735 ;
        RECT 73.650 179.480 73.910 179.800 ;
        RECT 73.710 174.360 73.850 179.480 ;
        RECT 75.030 179.140 75.290 179.460 ;
        RECT 75.090 177.760 75.230 179.140 ;
        RECT 76.515 177.925 78.055 178.295 ;
        RECT 75.030 177.440 75.290 177.760 ;
        RECT 79.230 175.040 79.370 185.600 ;
        RECT 79.815 180.645 81.355 181.015 ;
        RECT 81.470 176.760 81.730 177.080 ;
        RECT 79.815 175.205 81.355 175.575 ;
        RECT 79.170 174.720 79.430 175.040 ;
        RECT 73.650 174.040 73.910 174.360 ;
        RECT 81.530 174.020 81.670 176.760 ;
        RECT 75.490 173.700 75.750 174.020 ;
        RECT 81.470 173.700 81.730 174.020 ;
        RECT 75.550 172.320 75.690 173.700 ;
        RECT 76.515 172.485 78.055 172.855 ;
        RECT 75.490 172.000 75.750 172.320 ;
        RECT 81.530 171.640 81.670 173.700 ;
        RECT 75.030 171.320 75.290 171.640 ;
        RECT 81.470 171.320 81.730 171.640 ;
        RECT 75.090 166.880 75.230 171.320 ;
        RECT 81.470 170.300 81.730 170.620 ;
        RECT 79.815 169.765 81.355 170.135 ;
        RECT 81.530 169.000 81.670 170.300 ;
        RECT 81.070 168.860 81.670 169.000 ;
        RECT 76.515 167.045 78.055 167.415 ;
        RECT 75.030 166.560 75.290 166.880 ;
        RECT 81.070 165.860 81.210 168.860 ;
        RECT 81.470 165.880 81.730 166.200 ;
        RECT 81.010 165.540 81.270 165.860 ;
        RECT 76.870 164.860 77.130 165.180 ;
        RECT 76.930 163.140 77.070 164.860 ;
        RECT 79.815 164.325 81.355 164.695 ;
        RECT 75.490 162.820 75.750 163.140 ;
        RECT 76.870 162.820 77.130 163.140 ;
        RECT 79.170 162.820 79.430 163.140 ;
        RECT 7.395 148.055 8.255 158.425 ;
        RECT 75.550 155.320 75.690 162.820 ;
        RECT 76.515 161.605 78.055 161.975 ;
        RECT 79.230 157.020 79.370 162.820 ;
        RECT 79.815 158.885 81.355 159.255 ;
        RECT 79.170 156.700 79.430 157.020 ;
        RECT 76.515 156.165 78.055 156.535 ;
        RECT 75.490 155.000 75.750 155.320 ;
        RECT 75.030 154.320 75.290 154.640 ;
        RECT 75.090 153.280 75.230 154.320 ;
        RECT 79.815 153.445 81.355 153.815 ;
        RECT 75.030 152.960 75.290 153.280 ;
        RECT 81.530 152.260 81.670 165.880 ;
        RECT 81.470 151.940 81.730 152.260 ;
        RECT 76.515 150.725 78.055 151.095 ;
        RECT 81.990 150.560 82.130 186.710 ;
        RECT 83.830 185.920 83.970 187.300 ;
        RECT 84.290 187.280 84.430 189.340 ;
        RECT 84.230 186.960 84.490 187.280 ;
        RECT 85.150 186.620 85.410 186.940 ;
        RECT 83.770 185.600 84.030 185.920 ;
        RECT 85.210 185.240 85.350 186.620 ;
        RECT 85.150 184.920 85.410 185.240 ;
        RECT 87.050 184.560 87.190 189.340 ;
        RECT 87.970 184.900 88.110 190.020 ;
        RECT 93.890 189.340 94.150 189.660 ;
        RECT 94.350 189.340 94.610 189.660 ;
        RECT 88.590 188.805 90.130 189.175 ;
        RECT 93.950 187.960 94.090 189.340 ;
        RECT 94.410 188.640 94.550 189.340 ;
        RECT 94.350 188.320 94.610 188.640 ;
        RECT 93.890 187.640 94.150 187.960 ;
        RECT 89.290 186.960 89.550 187.280 ;
        RECT 89.350 185.920 89.490 186.960 ;
        RECT 91.890 186.085 93.430 186.455 ;
        RECT 89.290 185.600 89.550 185.920 ;
        RECT 94.410 185.240 94.550 188.320 ;
        RECT 94.870 187.620 95.010 190.020 ;
        RECT 100.390 189.400 100.530 190.360 ;
        RECT 99.930 189.260 100.530 189.400 ;
        RECT 99.930 188.720 100.070 189.260 ;
        RECT 100.665 188.805 102.205 189.175 ;
        RECT 99.930 188.580 100.530 188.720 ;
        RECT 94.810 187.300 95.070 187.620 ;
        RECT 99.870 187.300 100.130 187.620 ;
        RECT 98.490 186.960 98.750 187.280 ;
        RECT 98.550 185.920 98.690 186.960 ;
        RECT 98.490 185.600 98.750 185.920 ;
        RECT 98.950 185.600 99.210 185.920 ;
        RECT 99.930 185.680 100.070 187.300 ;
        RECT 94.350 184.920 94.610 185.240 ;
        RECT 87.910 184.580 88.170 184.900 ;
        RECT 91.130 184.580 91.390 184.900 ;
        RECT 86.990 184.240 87.250 184.560 ;
        RECT 83.770 183.900 84.030 184.220 ;
        RECT 83.830 183.200 83.970 183.900 ;
        RECT 87.970 183.200 88.110 184.580 ;
        RECT 88.590 183.365 90.130 183.735 ;
        RECT 91.190 183.200 91.330 184.580 ;
        RECT 92.970 184.240 93.230 184.560 ;
        RECT 83.770 182.880 84.030 183.200 ;
        RECT 87.910 182.880 88.170 183.200 ;
        RECT 91.130 182.880 91.390 183.200 ;
        RECT 93.030 182.180 93.170 184.240 ;
        RECT 94.410 183.200 94.550 184.920 ;
        RECT 95.730 183.900 95.990 184.220 ;
        RECT 94.350 182.880 94.610 183.200 ;
        RECT 95.790 182.180 95.930 183.900 ;
        RECT 99.010 182.860 99.150 185.600 ;
        RECT 99.470 185.540 100.070 185.680 ;
        RECT 98.950 182.540 99.210 182.860 ;
        RECT 92.970 181.860 93.230 182.180 ;
        RECT 95.730 181.860 95.990 182.180 ;
        RECT 93.890 181.520 94.150 181.840 ;
        RECT 91.890 180.645 93.430 181.015 ;
        RECT 82.390 179.480 82.650 179.800 ;
        RECT 82.450 174.360 82.590 179.480 ;
        RECT 85.610 178.800 85.870 179.120 ;
        RECT 85.150 178.460 85.410 178.780 ;
        RECT 85.210 177.080 85.350 178.460 ;
        RECT 85.150 176.760 85.410 177.080 ;
        RECT 82.850 176.420 83.110 176.740 ;
        RECT 82.390 174.040 82.650 174.360 ;
        RECT 82.910 173.760 83.050 176.420 ;
        RECT 83.770 176.080 84.030 176.400 ;
        RECT 82.450 173.620 83.050 173.760 ;
        RECT 82.450 171.640 82.590 173.620 ;
        RECT 82.850 173.020 83.110 173.340 ;
        RECT 82.390 171.320 82.650 171.640 ;
        RECT 82.450 168.580 82.590 171.320 ;
        RECT 82.910 171.300 83.050 173.020 ;
        RECT 83.830 172.320 83.970 176.080 ;
        RECT 83.770 172.000 84.030 172.320 ;
        RECT 82.850 170.980 83.110 171.300 ;
        RECT 83.830 168.580 83.970 172.000 ;
        RECT 85.670 168.920 85.810 178.800 ;
        RECT 88.590 177.925 90.130 178.295 ;
        RECT 91.890 175.205 93.430 175.575 ;
        RECT 93.950 174.360 94.090 181.520 ;
        RECT 99.470 180.480 99.610 185.540 ;
        RECT 100.390 184.900 100.530 188.580 ;
        RECT 101.250 186.960 101.510 187.280 ;
        RECT 101.310 185.240 101.450 186.960 ;
        RECT 102.690 186.940 102.830 192.400 ;
        RECT 106.770 192.060 107.030 192.380 ;
        RECT 103.965 191.525 105.505 191.895 ;
        RECT 106.310 191.040 106.570 191.360 ;
        RECT 103.090 190.360 103.350 190.680 ;
        RECT 104.470 190.360 104.730 190.680 ;
        RECT 102.630 186.620 102.890 186.940 ;
        RECT 102.690 185.240 102.830 186.620 ;
        RECT 103.150 185.240 103.290 190.360 ;
        RECT 104.010 190.020 104.270 190.340 ;
        RECT 103.550 189.340 103.810 189.660 ;
        RECT 103.610 185.920 103.750 189.340 ;
        RECT 104.070 188.640 104.210 190.020 ;
        RECT 104.010 188.320 104.270 188.640 ;
        RECT 104.530 187.960 104.670 190.360 ;
        RECT 106.370 188.300 106.510 191.040 ;
        RECT 106.310 187.980 106.570 188.300 ;
        RECT 104.470 187.640 104.730 187.960 ;
        RECT 103.965 186.085 105.505 186.455 ;
        RECT 106.370 185.920 106.510 187.980 ;
        RECT 106.830 187.620 106.970 192.060 ;
        RECT 111.430 191.360 111.570 192.400 ;
        RECT 116.040 191.525 117.580 191.895 ;
        RECT 111.370 191.040 111.630 191.360 ;
        RECT 107.690 190.700 107.950 191.020 ;
        RECT 107.750 188.640 107.890 190.700 ;
        RECT 109.070 190.360 109.330 190.680 ;
        RECT 107.690 188.320 107.950 188.640 ;
        RECT 108.150 187.640 108.410 187.960 ;
        RECT 106.770 187.300 107.030 187.620 ;
        RECT 103.550 185.600 103.810 185.920 ;
        RECT 106.310 185.600 106.570 185.920 ;
        RECT 101.250 184.920 101.510 185.240 ;
        RECT 102.630 184.920 102.890 185.240 ;
        RECT 103.090 184.920 103.350 185.240 ;
        RECT 100.330 184.580 100.590 184.900 ;
        RECT 100.390 183.960 100.530 184.580 ;
        RECT 99.930 183.820 100.530 183.960 ;
        RECT 99.930 183.280 100.070 183.820 ;
        RECT 100.665 183.365 102.205 183.735 ;
        RECT 99.930 183.140 100.530 183.280 ;
        RECT 100.390 181.500 100.530 183.140 ;
        RECT 102.630 181.520 102.890 181.840 ;
        RECT 100.330 181.180 100.590 181.500 ;
        RECT 99.410 180.160 99.670 180.480 ;
        RECT 99.870 179.820 100.130 180.140 ;
        RECT 97.110 178.460 97.370 178.780 ;
        RECT 96.190 177.100 96.450 177.420 ;
        RECT 93.890 174.040 94.150 174.360 ;
        RECT 93.430 173.020 93.690 173.340 ;
        RECT 88.590 172.485 90.130 172.855 ;
        RECT 93.490 171.640 93.630 173.020 ;
        RECT 93.430 171.320 93.690 171.640 ;
        RECT 86.530 170.640 86.790 170.960 ;
        RECT 85.610 168.600 85.870 168.920 ;
        RECT 82.390 168.260 82.650 168.580 ;
        RECT 83.770 168.260 84.030 168.580 ;
        RECT 82.450 166.200 82.590 168.260 ;
        RECT 82.390 165.880 82.650 166.200 ;
        RECT 85.610 165.540 85.870 165.860 ;
        RECT 85.670 164.160 85.810 165.540 ;
        RECT 85.610 163.840 85.870 164.160 ;
        RECT 82.850 162.140 83.110 162.460 ;
        RECT 84.230 162.140 84.490 162.460 ;
        RECT 82.910 158.380 83.050 162.140 ;
        RECT 84.290 161.440 84.430 162.140 ;
        RECT 84.230 161.120 84.490 161.440 ;
        RECT 82.850 158.060 83.110 158.380 ;
        RECT 82.390 157.720 82.650 158.040 ;
        RECT 82.450 156.000 82.590 157.720 ;
        RECT 82.390 155.680 82.650 156.000 ;
        RECT 82.910 154.980 83.050 158.060 ;
        RECT 85.610 157.380 85.870 157.700 ;
        RECT 82.850 154.660 83.110 154.980 ;
        RECT 84.230 154.660 84.490 154.980 ;
        RECT 82.910 151.920 83.050 154.660 ;
        RECT 82.850 151.600 83.110 151.920 ;
        RECT 84.290 151.580 84.430 154.660 ;
        RECT 84.690 153.980 84.950 154.300 ;
        RECT 84.750 153.280 84.890 153.980 ;
        RECT 84.690 152.960 84.950 153.280 ;
        RECT 84.230 151.260 84.490 151.580 ;
        RECT 81.930 150.240 82.190 150.560 ;
        RECT 20.350 149.765 20.770 150.185 ;
        RECT 84.290 149.880 84.430 151.260 ;
        RECT 84.230 149.560 84.490 149.880 ;
        RECT 81.930 149.220 82.190 149.540 ;
        RECT 14.840 148.055 16.515 148.550 ;
        RECT 7.395 147.645 16.515 148.055 ;
        RECT 7.395 109.610 8.255 147.645 ;
        RECT 14.840 147.275 16.515 147.645 ;
        RECT 19.600 147.505 20.050 147.925 ;
        RECT 49.000 147.760 50.500 148.755 ;
        RECT 79.815 148.005 81.355 148.375 ;
        RECT 21.010 142.895 21.425 143.355 ;
        RECT 25.335 143.245 26.440 144.355 ;
        RECT 80.610 141.660 81.210 141.800 ;
        RECT 80.610 141.310 80.750 141.660 ;
        RECT 19.810 140.425 24.780 140.705 ;
        RECT 18.925 139.415 19.155 139.430 ;
        RECT 18.885 139.350 19.205 139.415 ;
        RECT 18.885 139.155 20.895 139.350 ;
        RECT 18.925 139.120 20.895 139.155 ;
        RECT 18.925 139.115 19.155 139.120 ;
        RECT 20.665 136.390 20.895 139.120 ;
        RECT 20.665 136.160 21.595 136.390 ;
        RECT 21.365 135.585 21.595 136.160 ;
        RECT 24.500 135.665 24.780 140.425 ;
        RECT 80.540 140.035 80.820 141.310 ;
        RECT 81.070 141.120 81.210 141.660 ;
        RECT 81.990 141.120 82.130 149.220 ;
        RECT 85.670 149.200 85.810 157.380 ;
        RECT 86.060 154.720 86.340 154.835 ;
        RECT 86.590 154.720 86.730 170.640 ;
        RECT 91.890 169.765 93.430 170.135 ;
        RECT 93.950 168.920 94.090 174.040 ;
        RECT 96.250 174.020 96.390 177.100 ;
        RECT 97.170 176.740 97.310 178.460 ;
        RECT 99.930 177.760 100.070 179.820 ;
        RECT 100.390 179.800 100.530 181.180 ;
        RECT 100.330 179.480 100.590 179.800 ;
        RECT 100.665 177.925 102.205 178.295 ;
        RECT 99.870 177.440 100.130 177.760 ;
        RECT 97.110 176.420 97.370 176.740 ;
        RECT 96.650 176.080 96.910 176.400 ;
        RECT 96.190 173.700 96.450 174.020 ;
        RECT 96.710 170.620 96.850 176.080 ;
        RECT 97.170 174.360 97.310 176.420 ;
        RECT 99.930 175.040 100.070 177.440 ;
        RECT 99.870 174.720 100.130 175.040 ;
        RECT 97.110 174.040 97.370 174.360 ;
        RECT 100.665 172.485 102.205 172.855 ;
        RECT 96.650 170.300 96.910 170.620 ;
        RECT 90.210 168.600 90.470 168.920 ;
        RECT 93.890 168.600 94.150 168.920 ;
        RECT 88.590 167.045 90.130 167.415 ;
        RECT 90.270 165.180 90.410 168.600 ;
        RECT 93.890 167.580 94.150 167.900 ;
        RECT 94.810 167.580 95.070 167.900 ;
        RECT 95.730 167.580 95.990 167.900 ;
        RECT 93.950 165.600 94.090 167.580 ;
        RECT 94.870 166.200 95.010 167.580 ;
        RECT 94.810 165.880 95.070 166.200 ;
        RECT 93.950 165.460 94.550 165.600 ;
        RECT 89.290 164.860 89.550 165.180 ;
        RECT 90.210 164.860 90.470 165.180 ;
        RECT 93.890 164.860 94.150 165.180 ;
        RECT 89.350 164.160 89.490 164.860 ;
        RECT 89.290 163.840 89.550 164.160 ;
        RECT 88.590 161.605 90.130 161.975 ;
        RECT 87.910 159.420 88.170 159.740 ;
        RECT 87.970 157.700 88.110 159.420 ;
        RECT 87.910 157.380 88.170 157.700 ;
        RECT 90.270 157.360 90.410 164.860 ;
        RECT 91.890 164.325 93.430 164.695 ;
        RECT 93.950 162.460 94.090 164.860 ;
        RECT 94.410 163.820 94.550 165.460 ;
        RECT 95.790 165.180 95.930 167.580 ;
        RECT 95.730 164.860 95.990 165.180 ;
        RECT 95.790 164.160 95.930 164.860 ;
        RECT 95.730 163.840 95.990 164.160 ;
        RECT 94.350 163.500 94.610 163.820 ;
        RECT 93.890 162.140 94.150 162.460 ;
        RECT 91.890 158.885 93.430 159.255 ;
        RECT 93.430 157.720 93.690 158.040 ;
        RECT 90.210 157.040 90.470 157.360 ;
        RECT 88.590 156.165 90.130 156.535 ;
        RECT 86.060 154.580 86.730 154.720 ;
        RECT 93.490 154.720 93.630 157.720 ;
        RECT 93.950 155.320 94.090 162.140 ;
        RECT 95.790 158.380 95.930 163.840 ;
        RECT 95.730 158.060 95.990 158.380 ;
        RECT 94.350 156.700 94.610 157.020 ;
        RECT 94.410 156.000 94.550 156.700 ;
        RECT 94.350 155.680 94.610 156.000 ;
        RECT 93.890 155.000 94.150 155.320 ;
        RECT 93.490 154.580 94.090 154.720 ;
        RECT 95.790 154.640 95.930 158.060 ;
        RECT 86.060 154.465 86.340 154.580 ;
        RECT 93.950 154.300 94.090 154.580 ;
        RECT 95.730 154.320 95.990 154.640 ;
        RECT 93.890 153.980 94.150 154.300 ;
        RECT 91.890 153.445 93.430 153.815 ;
        RECT 93.950 152.260 94.090 153.980 ;
        RECT 96.710 152.940 96.850 170.300 ;
        RECT 100.665 167.045 102.205 167.415 ;
        RECT 100.665 161.605 102.205 161.975 ;
        RECT 102.690 161.100 102.830 181.520 ;
        RECT 103.150 177.760 103.290 184.920 ;
        RECT 106.310 184.640 106.570 184.900 ;
        RECT 106.830 184.640 106.970 187.300 ;
        RECT 108.210 185.920 108.350 187.640 ;
        RECT 108.150 185.600 108.410 185.920 ;
        RECT 106.310 184.580 106.970 184.640 ;
        RECT 106.370 184.500 106.970 184.580 ;
        RECT 105.850 181.520 106.110 181.840 ;
        RECT 103.965 180.645 105.505 181.015 ;
        RECT 105.910 179.800 106.050 181.520 ;
        RECT 106.370 181.500 106.510 184.500 ;
        RECT 106.770 183.900 107.030 184.220 ;
        RECT 106.310 181.180 106.570 181.500 ;
        RECT 105.850 179.480 106.110 179.800 ;
        RECT 103.090 177.440 103.350 177.760 ;
        RECT 103.550 176.420 103.810 176.740 ;
        RECT 103.610 175.040 103.750 176.420 ;
        RECT 105.850 175.740 106.110 176.060 ;
        RECT 103.965 175.205 105.505 175.575 ;
        RECT 103.550 174.720 103.810 175.040 ;
        RECT 103.090 170.640 103.350 170.960 ;
        RECT 103.150 169.600 103.290 170.640 ;
        RECT 103.965 169.765 105.505 170.135 ;
        RECT 105.910 169.600 106.050 175.740 ;
        RECT 106.370 174.700 106.510 181.180 ;
        RECT 106.830 179.800 106.970 183.900 ;
        RECT 107.690 180.160 107.950 180.480 ;
        RECT 106.770 179.480 107.030 179.800 ;
        RECT 107.230 175.740 107.490 176.060 ;
        RECT 107.290 175.040 107.430 175.740 ;
        RECT 107.230 174.720 107.490 175.040 ;
        RECT 106.310 174.380 106.570 174.700 ;
        RECT 107.750 174.360 107.890 180.160 ;
        RECT 108.610 176.420 108.870 176.740 ;
        RECT 108.670 175.040 108.810 176.420 ;
        RECT 108.610 174.720 108.870 175.040 ;
        RECT 107.690 174.040 107.950 174.360 ;
        RECT 103.090 169.280 103.350 169.600 ;
        RECT 105.850 169.280 106.110 169.600 ;
        RECT 107.750 168.920 107.890 174.040 ;
        RECT 108.610 173.700 108.870 174.020 ;
        RECT 108.670 172.320 108.810 173.700 ;
        RECT 108.610 172.000 108.870 172.320 ;
        RECT 108.150 170.300 108.410 170.620 ;
        RECT 107.690 168.600 107.950 168.920 ;
        RECT 108.210 167.900 108.350 170.300 ;
        RECT 108.150 167.580 108.410 167.900 ;
        RECT 106.310 166.560 106.570 166.880 ;
        RECT 103.965 164.325 105.505 164.695 ;
        RECT 106.370 161.440 106.510 166.560 ;
        RECT 106.770 164.860 107.030 165.180 ;
        RECT 106.310 161.120 106.570 161.440 ;
        RECT 102.630 160.780 102.890 161.100 ;
        RECT 102.170 160.100 102.430 160.420 ;
        RECT 102.230 158.720 102.370 160.100 ;
        RECT 102.170 158.400 102.430 158.720 ;
        RECT 102.690 157.360 102.830 160.780 ;
        RECT 103.090 160.100 103.350 160.420 ;
        RECT 103.150 158.040 103.290 160.100 ;
        RECT 103.550 159.420 103.810 159.740 ;
        RECT 103.090 157.720 103.350 158.040 ;
        RECT 102.630 157.040 102.890 157.360 ;
        RECT 100.665 156.165 102.205 156.535 ;
        RECT 102.170 153.980 102.430 154.300 ;
        RECT 102.230 152.940 102.370 153.980 ;
        RECT 96.650 152.620 96.910 152.940 ;
        RECT 102.170 152.620 102.430 152.940 ;
        RECT 93.890 151.940 94.150 152.260 ;
        RECT 86.070 151.600 86.330 151.920 ;
        RECT 86.130 151.180 86.270 151.600 ;
        RECT 86.130 151.040 87.650 151.180 ;
        RECT 87.510 149.200 87.650 151.040 ;
        RECT 88.590 150.725 90.130 151.095 ;
        RECT 93.950 150.560 94.090 151.940 ;
        RECT 102.690 151.920 102.830 157.040 ;
        RECT 103.090 156.700 103.350 157.020 ;
        RECT 103.150 156.000 103.290 156.700 ;
        RECT 103.090 155.680 103.350 156.000 ;
        RECT 103.610 154.640 103.750 159.420 ;
        RECT 103.965 158.885 105.505 159.255 ;
        RECT 104.930 157.440 105.190 157.700 ;
        RECT 106.370 157.440 106.510 161.120 ;
        RECT 104.930 157.380 106.510 157.440 ;
        RECT 104.990 157.300 106.510 157.380 ;
        RECT 104.470 156.700 104.730 157.020 ;
        RECT 104.530 156.000 104.670 156.700 ;
        RECT 106.830 156.080 106.970 164.860 ;
        RECT 108.210 163.140 108.350 167.580 ;
        RECT 108.150 162.820 108.410 163.140 ;
        RECT 104.470 155.680 104.730 156.000 ;
        RECT 106.830 155.940 107.430 156.080 ;
        RECT 106.770 155.340 107.030 155.660 ;
        RECT 103.550 154.320 103.810 154.640 ;
        RECT 103.090 153.980 103.350 154.300 ;
        RECT 103.150 152.600 103.290 153.980 ;
        RECT 103.965 153.445 105.505 153.815 ;
        RECT 103.090 152.280 103.350 152.600 ;
        RECT 105.390 152.280 105.650 152.600 ;
        RECT 102.630 151.600 102.890 151.920 ;
        RECT 100.665 150.725 102.205 151.095 ;
        RECT 102.690 150.560 102.830 151.600 ;
        RECT 105.450 150.560 105.590 152.280 ;
        RECT 93.890 150.240 94.150 150.560 ;
        RECT 102.630 150.240 102.890 150.560 ;
        RECT 105.390 150.240 105.650 150.560 ;
        RECT 106.830 149.540 106.970 155.340 ;
        RECT 107.290 153.280 107.430 155.940 ;
        RECT 108.210 155.320 108.350 162.820 ;
        RECT 108.610 160.100 108.870 160.420 ;
        RECT 108.670 157.700 108.810 160.100 ;
        RECT 108.610 157.380 108.870 157.700 ;
        RECT 108.670 156.000 108.810 157.380 ;
        RECT 108.610 155.680 108.870 156.000 ;
        RECT 108.150 155.000 108.410 155.320 ;
        RECT 107.230 152.960 107.490 153.280 ;
        RECT 107.290 150.220 107.430 152.960 ;
        RECT 107.230 149.900 107.490 150.220 ;
        RECT 106.770 149.220 107.030 149.540 ;
        RECT 85.610 148.880 85.870 149.200 ;
        RECT 87.450 148.880 87.710 149.200 ;
        RECT 109.130 148.860 109.270 190.360 ;
        RECT 120.110 189.680 120.370 190.000 ;
        RECT 111.830 189.340 112.090 189.660 ;
        RECT 120.170 189.515 120.310 189.680 ;
        RECT 111.890 187.960 112.030 189.340 ;
        RECT 112.740 188.805 114.280 189.175 ;
        RECT 120.100 189.145 120.380 189.515 ;
        RECT 119.190 188.320 119.450 188.640 ;
        RECT 111.830 187.640 112.090 187.960 ;
        RECT 113.210 186.620 113.470 186.940 ;
        RECT 113.270 185.580 113.410 186.620 ;
        RECT 116.040 186.085 117.580 186.455 ;
        RECT 113.210 185.260 113.470 185.580 ;
        RECT 110.910 184.580 111.170 184.900 ;
        RECT 110.970 180.480 111.110 184.580 ;
        RECT 112.740 183.365 114.280 183.735 ;
        RECT 115.050 181.520 115.310 181.840 ;
        RECT 111.830 181.180 112.090 181.500 ;
        RECT 110.910 180.160 111.170 180.480 ;
        RECT 111.370 176.760 111.630 177.080 ;
        RECT 111.430 174.020 111.570 176.760 ;
        RECT 111.890 175.040 112.030 181.180 ;
        RECT 112.290 178.460 112.550 178.780 ;
        RECT 112.350 176.740 112.490 178.460 ;
        RECT 112.740 177.925 114.280 178.295 ;
        RECT 115.110 177.760 115.250 181.520 ;
        RECT 116.040 180.645 117.580 181.015 ;
        RECT 115.050 177.440 115.310 177.760 ;
        RECT 118.730 176.760 118.990 177.080 ;
        RECT 112.290 176.420 112.550 176.740 ;
        RECT 114.590 175.740 114.850 176.060 ;
        RECT 115.050 175.740 115.310 176.060 ;
        RECT 115.510 175.740 115.770 176.060 ;
        RECT 117.810 175.740 118.070 176.060 ;
        RECT 111.830 174.720 112.090 175.040 ;
        RECT 111.370 173.700 111.630 174.020 ;
        RECT 112.740 172.485 114.280 172.855 ;
        RECT 114.130 170.300 114.390 170.620 ;
        RECT 114.190 169.600 114.330 170.300 ;
        RECT 114.130 169.280 114.390 169.600 ;
        RECT 112.740 167.045 114.280 167.415 ;
        RECT 114.650 166.280 114.790 175.740 ;
        RECT 115.110 174.020 115.250 175.740 ;
        RECT 115.050 173.700 115.310 174.020 ;
        RECT 115.050 173.020 115.310 173.340 ;
        RECT 115.110 171.640 115.250 173.020 ;
        RECT 115.050 171.320 115.310 171.640 ;
        RECT 115.570 166.880 115.710 175.740 ;
        RECT 116.040 175.205 117.580 175.575 ;
        RECT 117.870 174.360 118.010 175.740 ;
        RECT 117.350 174.040 117.610 174.360 ;
        RECT 117.810 174.040 118.070 174.360 ;
        RECT 117.410 171.980 117.550 174.040 ;
        RECT 117.350 171.660 117.610 171.980 ;
        RECT 116.040 169.765 117.580 170.135 ;
        RECT 117.870 169.600 118.010 174.040 ;
        RECT 118.270 173.020 118.530 173.340 ;
        RECT 117.810 169.280 118.070 169.600 ;
        RECT 115.510 166.560 115.770 166.880 ;
        RECT 114.650 166.140 115.250 166.280 ;
        RECT 114.590 165.540 114.850 165.860 ;
        RECT 110.450 164.860 110.710 165.180 ;
        RECT 111.830 164.860 112.090 165.180 ;
        RECT 109.530 162.140 109.790 162.460 ;
        RECT 109.590 160.420 109.730 162.140 ;
        RECT 110.510 160.420 110.650 164.860 ;
        RECT 111.890 163.820 112.030 164.860 ;
        RECT 111.830 163.500 112.090 163.820 ;
        RECT 112.740 161.605 114.280 161.975 ;
        RECT 114.650 161.440 114.790 165.540 ;
        RECT 115.110 165.180 115.250 166.140 ;
        RECT 118.330 165.520 118.470 173.020 ;
        RECT 118.270 165.200 118.530 165.520 ;
        RECT 115.050 164.860 115.310 165.180 ;
        RECT 116.040 164.325 117.580 164.695 ;
        RECT 115.050 162.140 115.310 162.460 ;
        RECT 114.590 161.120 114.850 161.440 ;
        RECT 115.110 160.760 115.250 162.140 ;
        RECT 115.050 160.440 115.310 160.760 ;
        RECT 109.530 160.100 109.790 160.420 ;
        RECT 110.450 160.100 110.710 160.420 ;
        RECT 109.590 158.040 109.730 160.100 ;
        RECT 109.530 157.720 109.790 158.040 ;
        RECT 109.590 154.980 109.730 157.720 ;
        RECT 110.510 157.020 110.650 160.100 ;
        RECT 115.110 158.040 115.250 160.440 ;
        RECT 116.040 158.885 117.580 159.255 ;
        RECT 118.790 158.040 118.930 176.760 ;
        RECT 115.050 157.720 115.310 158.040 ;
        RECT 118.730 157.720 118.990 158.040 ;
        RECT 110.910 157.380 111.170 157.700 ;
        RECT 115.510 157.380 115.770 157.700 ;
        RECT 110.450 156.700 110.710 157.020 ;
        RECT 109.530 154.660 109.790 154.980 ;
        RECT 110.970 153.280 111.110 157.380 ;
        RECT 112.740 156.165 114.280 156.535 ;
        RECT 115.570 156.000 115.710 157.380 ;
        RECT 115.510 155.680 115.770 156.000 ;
        RECT 117.810 155.680 118.070 156.000 ;
        RECT 115.050 154.320 115.310 154.640 ;
        RECT 115.110 153.280 115.250 154.320 ;
        RECT 116.040 153.445 117.580 153.815 ;
        RECT 110.910 152.960 111.170 153.280 ;
        RECT 115.050 152.960 115.310 153.280 ;
        RECT 110.970 149.880 111.110 152.960 ;
        RECT 114.590 151.260 114.850 151.580 ;
        RECT 112.740 150.725 114.280 151.095 ;
        RECT 114.650 150.560 114.790 151.260 ;
        RECT 114.590 150.240 114.850 150.560 ;
        RECT 117.870 149.880 118.010 155.680 ;
        RECT 119.250 153.280 119.390 188.320 ;
        RECT 120.100 153.785 120.380 154.155 ;
        RECT 120.170 153.280 120.310 153.785 ;
        RECT 119.190 152.960 119.450 153.280 ;
        RECT 120.110 152.960 120.370 153.280 ;
        RECT 110.910 149.560 111.170 149.880 ;
        RECT 117.810 149.560 118.070 149.880 ;
        RECT 109.530 148.880 109.790 149.200 ;
        RECT 109.070 148.540 109.330 148.860 ;
        RECT 91.890 148.005 93.430 148.375 ;
        RECT 103.965 148.005 105.505 148.375 ;
        RECT 109.590 143.840 109.730 148.880 ;
        RECT 116.040 148.005 117.580 148.375 ;
        RECT 109.590 143.700 110.650 143.840 ;
        RECT 110.510 141.310 110.650 143.700 ;
        RECT 81.070 140.980 82.130 141.120 ;
        RECT 80.195 138.950 81.260 140.035 ;
        RECT 110.440 139.950 110.720 141.310 ;
        RECT 110.180 139.050 111.080 139.950 ;
        RECT 80.540 137.310 80.820 138.950 ;
        RECT 110.440 137.310 110.720 139.050 ;
        RECT 88.130 135.875 152.705 135.900 ;
        RECT 21.350 135.265 21.610 135.585 ;
        RECT 24.470 135.385 24.810 135.665 ;
        RECT 88.110 135.325 152.705 135.875 ;
        RECT 88.130 135.300 152.705 135.325 ;
        RECT 21.950 133.825 22.340 134.145 ;
        RECT 24.010 133.855 24.340 134.135 ;
        RECT 22.020 133.705 22.240 133.825 ;
        RECT 17.500 131.110 18.040 131.560 ;
        RECT 19.640 131.270 19.900 131.365 ;
        RECT 22.045 131.270 22.195 133.705 ;
        RECT 19.640 131.120 22.195 131.270 ;
        RECT 12.350 123.435 14.535 125.235 ;
        RECT 17.620 121.155 17.910 131.110 ;
        RECT 19.640 131.045 19.900 131.120 ;
        RECT 24.100 130.775 24.260 133.855 ;
        RECT 23.910 130.405 24.310 130.775 ;
        RECT 46.315 121.625 47.120 122.425 ;
        RECT 46.570 121.155 46.860 121.625 ;
        RECT 17.620 120.865 103.915 121.155 ;
        RECT 20.130 111.795 20.550 112.215 ;
        RECT 14.230 109.610 15.745 109.985 ;
        RECT 7.395 109.085 15.745 109.610 ;
        RECT 19.380 109.535 19.830 109.955 ;
        RECT 103.625 109.320 103.915 120.865 ;
        RECT 1.000 82.525 2.500 83.410 ;
        RECT 7.395 73.120 8.255 109.085 ;
        RECT 14.230 108.720 15.745 109.085 ;
        RECT 103.490 108.900 104.040 109.320 ;
        RECT 72.460 107.210 139.730 107.470 ;
        RECT 20.790 104.925 21.205 105.385 ;
        RECT 25.115 105.275 26.220 106.385 ;
        RECT 19.590 102.455 24.560 102.735 ;
        RECT 18.705 101.445 18.935 101.460 ;
        RECT 18.665 101.380 18.985 101.445 ;
        RECT 18.665 101.185 20.675 101.380 ;
        RECT 18.705 101.150 20.675 101.185 ;
        RECT 18.705 101.145 18.935 101.150 ;
        RECT 20.445 98.420 20.675 101.150 ;
        RECT 20.445 98.190 21.375 98.420 ;
        RECT 21.145 97.615 21.375 98.190 ;
        RECT 24.280 97.695 24.560 102.455 ;
        RECT 21.130 97.295 21.390 97.615 ;
        RECT 24.250 97.415 24.590 97.695 ;
        RECT 21.730 95.855 22.120 96.175 ;
        RECT 23.790 95.885 24.120 96.165 ;
        RECT 21.800 95.735 22.020 95.855 ;
        RECT 19.420 93.300 19.680 93.395 ;
        RECT 21.825 93.300 21.975 95.735 ;
        RECT 19.420 93.150 21.975 93.300 ;
        RECT 19.420 93.120 19.680 93.150 ;
        RECT 19.410 93.075 19.680 93.120 ;
        RECT 19.410 85.070 19.670 93.075 ;
        RECT 23.880 92.805 24.040 95.885 ;
        RECT 23.690 92.435 24.090 92.805 ;
        RECT 44.310 88.715 45.115 89.515 ;
        RECT 44.605 85.070 44.865 88.715 ;
        RECT 49.000 88.350 50.500 89.630 ;
        RECT 72.460 85.070 72.720 107.210 ;
        RECT 19.410 84.810 72.720 85.070 ;
        RECT 42.625 76.380 43.490 79.340 ;
        RECT 42.615 75.545 43.490 76.380 ;
        RECT 7.390 72.580 8.255 73.120 ;
        RECT 42.625 74.150 43.490 75.545 ;
        RECT 42.625 73.115 43.500 74.150 ;
        RECT 1.000 63.980 2.500 64.120 ;
        RECT 7.395 63.980 8.255 72.580 ;
        RECT 1.000 62.700 8.255 63.980 ;
        RECT 1.000 62.600 2.500 62.700 ;
        RECT 7.395 56.030 8.255 62.700 ;
        RECT 14.580 72.450 23.770 72.710 ;
        RECT 14.580 49.390 14.840 72.450 ;
        RECT 23.510 72.300 23.770 72.450 ;
        RECT 23.400 71.850 23.830 72.300 ;
        RECT 32.795 71.800 33.470 72.475 ;
        RECT 27.400 69.580 28.085 70.140 ;
        RECT 42.625 69.770 43.490 73.115 ;
        RECT 48.990 69.770 50.510 70.220 ;
        RECT 42.625 68.650 50.510 69.770 ;
        RECT 27.310 67.270 27.900 67.900 ;
        RECT 35.135 65.930 35.590 65.975 ;
        RECT 42.625 65.930 43.490 68.650 ;
        RECT 48.990 68.440 50.510 68.650 ;
        RECT 35.135 65.670 43.490 65.930 ;
        RECT 35.135 65.595 35.590 65.670 ;
        RECT 34.430 64.585 34.980 65.080 ;
        RECT 34.455 64.580 34.835 64.585 ;
        RECT 18.930 63.285 19.550 63.720 ;
        RECT 19.070 60.435 19.415 63.285 ;
        RECT 27.550 63.225 28.240 63.780 ;
        RECT 42.625 60.435 43.490 65.670 ;
        RECT 53.130 61.095 54.030 61.775 ;
        RECT 19.070 60.090 43.490 60.435 ;
        RECT 28.685 59.095 29.310 59.605 ;
        RECT 28.690 59.090 29.305 59.095 ;
        RECT 33.990 59.080 34.890 59.725 ;
        RECT 26.380 58.435 27.145 58.735 ;
        RECT 26.380 58.040 29.665 58.435 ;
        RECT 26.380 57.705 27.145 58.040 ;
        RECT 22.730 56.360 23.980 57.440 ;
        RECT 23.060 49.390 25.760 50.500 ;
        RECT 14.580 49.130 25.760 49.390 ;
        RECT 23.060 48.560 25.760 49.130 ;
        RECT 0.995 35.135 2.505 36.290 ;
        RECT 7.855 29.580 8.595 29.690 ;
        RECT 28.975 29.580 29.665 58.040 ;
        RECT 42.625 56.030 43.490 60.090 ;
        RECT 55.390 56.715 56.290 57.505 ;
        RECT 88.130 39.290 88.730 102.460 ;
        RECT 103.270 101.850 104.190 102.460 ;
        RECT 103.570 97.225 103.850 101.850 ;
        RECT 139.450 97.225 139.730 107.210 ;
        RECT 101.235 88.755 102.775 89.125 ;
        RECT 103.640 88.590 103.780 97.225 ;
        RECT 116.530 88.755 118.070 89.125 ;
        RECT 131.825 88.755 133.365 89.125 ;
        RECT 139.520 88.590 139.660 97.225 ;
        RECT 147.120 88.755 148.660 89.125 ;
        RECT 151.870 89.095 152.150 89.465 ;
        RECT 103.580 88.270 103.840 88.590 ;
        RECT 139.460 88.270 139.720 88.590 ;
        RECT 151.940 88.250 152.080 89.095 ;
        RECT 151.880 87.930 152.140 88.250 ;
        RECT 106.340 87.590 106.600 87.910 ;
        RECT 140.380 87.590 140.640 87.910 ;
        RECT 97.935 86.035 99.475 86.405 ;
        RECT 101.235 83.315 102.775 83.685 ;
        RECT 97.935 80.595 99.475 80.965 ;
        RECT 105.870 79.575 106.150 79.945 ;
        RECT 101.235 77.875 102.775 78.245 ;
        RECT 97.935 75.155 99.475 75.525 ;
        RECT 105.940 74.990 106.080 79.575 ;
        RECT 105.880 74.670 106.140 74.990 ;
        RECT 101.235 72.435 102.775 72.805 ;
        RECT 97.935 69.715 99.475 70.085 ;
        RECT 103.580 68.210 103.840 68.530 ;
        RECT 100.360 67.530 100.620 67.850 ;
        RECT 100.420 66.490 100.560 67.530 ;
        RECT 101.235 66.995 102.775 67.365 ;
        RECT 100.360 66.170 100.620 66.490 ;
        RECT 101.740 64.810 102.000 65.130 ;
        RECT 103.120 64.810 103.380 65.130 ;
        RECT 97.935 64.275 99.475 64.645 ;
        RECT 101.800 64.110 101.940 64.810 ;
        RECT 101.740 63.790 102.000 64.110 ;
        RECT 100.360 62.430 100.620 62.750 ;
        RECT 93.000 62.090 93.260 62.410 ;
        RECT 93.060 61.390 93.200 62.090 ;
        RECT 100.420 61.390 100.560 62.430 ;
        RECT 103.180 62.410 103.320 64.810 ;
        RECT 103.120 62.090 103.380 62.410 ;
        RECT 101.235 61.555 102.775 61.925 ;
        RECT 93.000 61.070 93.260 61.390 ;
        RECT 95.760 61.070 96.020 61.390 ;
        RECT 100.360 61.070 100.620 61.390 ;
        RECT 92.540 51.890 92.800 52.210 ;
        RECT 92.600 50.170 92.740 51.890 ;
        RECT 92.540 49.850 92.800 50.170 ;
        RECT 92.600 47.790 92.740 49.850 ;
        RECT 92.540 47.470 92.800 47.790 ;
        RECT 90.240 41.010 90.500 41.330 ;
        RECT 88.105 38.625 88.790 39.290 ;
        RECT 90.300 39.145 90.440 41.010 ;
        RECT 90.230 38.775 90.510 39.145 ;
        RECT 95.820 38.610 95.960 61.070 ;
        RECT 98.060 60.390 98.320 60.710 ;
        RECT 99.440 60.390 99.700 60.710 ;
        RECT 99.900 60.390 100.160 60.710 ;
        RECT 102.200 60.390 102.460 60.710 ;
        RECT 98.120 59.940 98.260 60.390 ;
        RECT 97.200 59.800 98.260 59.940 ;
        RECT 96.680 59.370 96.940 59.690 ;
        RECT 96.740 58.670 96.880 59.370 ;
        RECT 96.680 58.350 96.940 58.670 ;
        RECT 97.200 57.310 97.340 59.800 ;
        RECT 99.500 59.690 99.640 60.390 ;
        RECT 99.440 59.370 99.700 59.690 ;
        RECT 97.935 58.835 99.475 59.205 ;
        RECT 99.960 58.670 100.100 60.390 ;
        RECT 100.820 60.050 101.080 60.370 ;
        RECT 100.880 58.670 101.020 60.050 ;
        RECT 99.900 58.350 100.160 58.670 ;
        RECT 100.820 58.350 101.080 58.670 ;
        RECT 102.260 57.650 102.400 60.390 ;
        RECT 97.600 57.330 97.860 57.650 ;
        RECT 98.980 57.330 99.240 57.650 ;
        RECT 100.360 57.330 100.620 57.650 ;
        RECT 102.200 57.330 102.460 57.650 ;
        RECT 97.140 56.990 97.400 57.310 ;
        RECT 96.680 56.650 96.940 56.970 ;
        RECT 96.740 53.230 96.880 56.650 ;
        RECT 97.660 55.950 97.800 57.330 ;
        RECT 97.600 55.630 97.860 55.950 ;
        RECT 99.040 55.270 99.180 57.330 ;
        RECT 100.420 55.270 100.560 57.330 ;
        RECT 101.235 56.115 102.775 56.485 ;
        RECT 103.180 55.270 103.320 62.090 ;
        RECT 103.640 61.390 103.780 68.210 ;
        RECT 105.880 62.090 106.140 62.410 ;
        RECT 103.580 61.070 103.840 61.390 ;
        RECT 104.960 60.390 105.220 60.710 ;
        RECT 98.980 54.950 99.240 55.270 ;
        RECT 100.360 54.950 100.620 55.270 ;
        RECT 103.120 54.950 103.380 55.270 ;
        RECT 97.935 53.395 99.475 53.765 ;
        RECT 96.680 52.910 96.940 53.230 ;
        RECT 100.420 51.530 100.560 54.950 ;
        RECT 103.180 52.210 103.320 54.950 ;
        RECT 100.820 51.890 101.080 52.210 ;
        RECT 103.120 51.890 103.380 52.210 ;
        RECT 100.360 51.210 100.620 51.530 ;
        RECT 97.140 49.170 97.400 49.490 ;
        RECT 96.220 48.490 96.480 48.810 ;
        RECT 96.280 47.110 96.420 48.490 ;
        RECT 96.220 46.790 96.480 47.110 ;
        RECT 97.200 44.730 97.340 49.170 ;
        RECT 99.900 48.490 100.160 48.810 ;
        RECT 97.935 47.955 99.475 48.325 ;
        RECT 99.960 46.770 100.100 48.490 ;
        RECT 99.900 46.450 100.160 46.770 ;
        RECT 97.140 44.410 97.400 44.730 ;
        RECT 96.220 43.050 96.480 43.370 ;
        RECT 96.280 40.650 96.420 43.050 ;
        RECT 97.935 42.515 99.475 42.885 ;
        RECT 96.220 40.330 96.480 40.650 ;
        RECT 95.760 38.290 96.020 38.610 ;
        RECT 96.680 38.290 96.940 38.610 ;
        RECT 98.980 38.465 99.240 38.610 ;
        RECT 95.820 36.230 95.960 38.290 ;
        RECT 96.740 36.570 96.880 38.290 ;
        RECT 98.970 38.095 99.250 38.465 ;
        RECT 99.900 37.610 100.160 37.930 ;
        RECT 100.420 37.670 100.560 51.210 ;
        RECT 100.880 50.420 101.020 51.890 ;
        RECT 104.040 51.550 104.300 51.870 ;
        RECT 101.235 50.675 102.775 51.045 ;
        RECT 100.880 50.280 101.480 50.420 ;
        RECT 101.340 49.830 101.480 50.280 ;
        RECT 101.280 49.510 101.540 49.830 ;
        RECT 104.100 49.490 104.240 51.550 ;
        RECT 100.820 49.170 101.080 49.490 ;
        RECT 104.040 49.170 104.300 49.490 ;
        RECT 100.880 45.070 101.020 49.170 ;
        RECT 101.235 45.235 102.775 45.605 ;
        RECT 100.820 44.750 101.080 45.070 ;
        RECT 104.100 44.390 104.240 49.170 ;
        RECT 104.040 44.070 104.300 44.390 ;
        RECT 101.235 39.795 102.775 40.165 ;
        RECT 102.200 39.310 102.460 39.630 ;
        RECT 100.820 37.950 101.080 38.270 ;
        RECT 100.880 37.670 101.020 37.950 ;
        RECT 97.935 37.075 99.475 37.445 ;
        RECT 99.960 36.910 100.100 37.610 ;
        RECT 100.420 37.530 101.020 37.670 ;
        RECT 99.900 36.590 100.160 36.910 ;
        RECT 96.680 36.250 96.940 36.570 ;
        RECT 100.420 36.230 100.560 37.530 ;
        RECT 102.260 36.570 102.400 39.310 ;
        RECT 104.040 38.290 104.300 38.610 ;
        RECT 103.580 37.950 103.840 38.270 ;
        RECT 102.200 36.250 102.460 36.570 ;
        RECT 95.760 35.910 96.020 36.230 ;
        RECT 100.360 35.910 100.620 36.230 ;
        RECT 93.460 35.570 93.720 35.890 ;
        RECT 93.520 31.470 93.660 35.570 ;
        RECT 95.820 35.210 95.960 35.910 ;
        RECT 103.640 35.890 103.780 37.950 ;
        RECT 100.820 35.570 101.080 35.890 ;
        RECT 103.580 35.570 103.840 35.890 ;
        RECT 95.760 34.890 96.020 35.210 ;
        RECT 99.900 34.890 100.160 35.210 ;
        RECT 99.960 34.190 100.100 34.890 ;
        RECT 100.880 34.190 101.020 35.570 ;
        RECT 101.235 34.355 102.775 34.725 ;
        RECT 99.900 33.870 100.160 34.190 ;
        RECT 100.820 33.870 101.080 34.190 ;
        RECT 102.200 33.870 102.460 34.190 ;
        RECT 99.900 33.190 100.160 33.510 ;
        RECT 97.935 31.635 99.475 32.005 ;
        RECT 99.960 31.470 100.100 33.190 ;
        RECT 102.260 32.490 102.400 33.870 ;
        RECT 103.640 33.590 103.780 35.570 ;
        RECT 102.720 33.510 103.780 33.590 ;
        RECT 104.100 33.510 104.240 38.290 ;
        RECT 105.020 37.930 105.160 60.390 ;
        RECT 105.940 60.030 106.080 62.090 ;
        RECT 105.880 59.710 106.140 60.030 ;
        RECT 105.940 49.490 106.080 59.710 ;
        RECT 106.400 52.550 106.540 87.590 ;
        RECT 113.230 86.035 114.770 86.405 ;
        RECT 128.525 86.035 130.065 86.405 ;
        RECT 118.300 84.870 118.560 85.190 ;
        RECT 125.660 84.870 125.920 85.190 ;
        RECT 116.530 83.315 118.070 83.685 ;
        RECT 118.360 82.130 118.500 84.870 ;
        RECT 121.980 84.530 122.240 84.850 ;
        RECT 122.440 84.530 122.700 84.850 ;
        RECT 122.040 82.810 122.180 84.530 ;
        RECT 122.500 83.150 122.640 84.530 ;
        RECT 122.900 83.850 123.160 84.170 ;
        RECT 124.740 83.850 125.000 84.170 ;
        RECT 122.440 82.830 122.700 83.150 ;
        RECT 118.760 82.490 119.020 82.810 ;
        RECT 121.980 82.490 122.240 82.810 ;
        RECT 113.240 81.810 113.500 82.130 ;
        RECT 115.080 81.810 115.340 82.130 ;
        RECT 118.300 81.810 118.560 82.130 ;
        RECT 113.300 81.360 113.440 81.810 ;
        RECT 112.840 81.220 113.440 81.360 ;
        RECT 112.840 80.390 112.980 81.220 ;
        RECT 113.230 80.595 114.770 80.965 ;
        RECT 112.840 80.250 113.440 80.390 ;
        RECT 110.940 79.430 111.200 79.750 ;
        RECT 107.260 75.690 107.520 76.010 ;
        RECT 107.320 73.630 107.460 75.690 ;
        RECT 111.000 73.970 111.140 79.430 ;
        RECT 113.300 76.690 113.440 80.250 ;
        RECT 115.140 79.070 115.280 81.810 ;
        RECT 115.540 81.130 115.800 81.450 ;
        RECT 115.080 78.750 115.340 79.070 ;
        RECT 115.600 78.730 115.740 81.130 ;
        RECT 118.360 79.750 118.500 81.810 ;
        RECT 118.300 79.430 118.560 79.750 ;
        RECT 115.540 78.410 115.800 78.730 ;
        RECT 116.530 77.875 118.070 78.245 ;
        RECT 115.080 76.710 115.340 77.030 ;
        RECT 118.300 76.710 118.560 77.030 ;
        RECT 113.240 76.430 113.500 76.690 ;
        RECT 112.840 76.370 113.500 76.430 ;
        RECT 112.840 76.290 113.440 76.370 ;
        RECT 110.940 73.650 111.200 73.970 ;
        RECT 107.260 73.310 107.520 73.630 ;
        RECT 109.100 73.310 109.360 73.630 ;
        RECT 109.160 72.270 109.300 73.310 ;
        RECT 109.100 71.950 109.360 72.270 ;
        RECT 109.560 71.270 109.820 71.590 ;
        RECT 109.620 66.830 109.760 71.270 ;
        RECT 111.000 68.870 111.140 73.650 ;
        RECT 112.840 71.590 112.980 76.290 ;
        RECT 113.230 75.155 114.770 75.525 ;
        RECT 115.140 72.270 115.280 76.710 ;
        RECT 115.540 74.670 115.800 74.990 ;
        RECT 115.080 71.950 115.340 72.270 ;
        RECT 112.780 71.270 113.040 71.590 ;
        RECT 115.080 70.250 115.340 70.570 ;
        RECT 113.230 69.715 114.770 70.085 ;
        RECT 115.140 68.870 115.280 70.250 ;
        RECT 110.940 68.550 111.200 68.870 ;
        RECT 115.080 68.550 115.340 68.870 ;
        RECT 109.560 66.510 109.820 66.830 ;
        RECT 107.260 64.810 107.520 65.130 ;
        RECT 107.320 63.430 107.460 64.810 ;
        RECT 107.260 63.340 107.520 63.430 ;
        RECT 106.860 63.200 107.520 63.340 ;
        RECT 106.860 60.710 107.000 63.200 ;
        RECT 107.260 63.110 107.520 63.200 ;
        RECT 107.260 62.090 107.520 62.410 ;
        RECT 107.720 62.090 107.980 62.410 ;
        RECT 107.320 61.390 107.460 62.090 ;
        RECT 107.260 61.070 107.520 61.390 ;
        RECT 107.780 60.790 107.920 62.090 ;
        RECT 107.320 60.710 107.920 60.790 ;
        RECT 106.800 60.390 107.060 60.710 ;
        RECT 107.260 60.650 107.920 60.710 ;
        RECT 107.260 60.390 107.520 60.650 ;
        RECT 107.320 58.670 107.460 60.390 ;
        RECT 108.640 59.370 108.900 59.690 ;
        RECT 107.260 58.350 107.520 58.670 ;
        RECT 108.700 54.250 108.840 59.370 ;
        RECT 108.640 53.930 108.900 54.250 ;
        RECT 106.340 52.230 106.600 52.550 ;
        RECT 106.800 51.550 107.060 51.870 ;
        RECT 107.720 51.550 107.980 51.870 ;
        RECT 106.860 50.170 107.000 51.550 ;
        RECT 107.780 50.510 107.920 51.550 ;
        RECT 108.180 51.210 108.440 51.530 ;
        RECT 107.720 50.190 107.980 50.510 ;
        RECT 106.800 49.850 107.060 50.170 ;
        RECT 106.860 49.490 107.000 49.850 ;
        RECT 105.880 49.170 106.140 49.490 ;
        RECT 106.800 49.170 107.060 49.490 ;
        RECT 105.420 48.490 105.680 48.810 ;
        RECT 105.480 46.090 105.620 48.490 ;
        RECT 105.420 45.770 105.680 46.090 ;
        RECT 105.480 44.390 105.620 45.770 ;
        RECT 105.940 44.730 106.080 49.170 ;
        RECT 107.780 47.790 107.920 50.190 ;
        RECT 108.240 47.790 108.380 51.210 ;
        RECT 107.260 47.470 107.520 47.790 ;
        RECT 107.720 47.470 107.980 47.790 ;
        RECT 108.180 47.470 108.440 47.790 ;
        RECT 107.320 47.190 107.460 47.470 ;
        RECT 108.700 47.190 108.840 53.930 ;
        RECT 109.100 51.210 109.360 51.530 ;
        RECT 109.160 50.510 109.300 51.210 ;
        RECT 109.100 50.190 109.360 50.510 ;
        RECT 107.320 47.050 108.840 47.190 ;
        RECT 105.880 44.410 106.140 44.730 ;
        RECT 105.420 44.070 105.680 44.390 ;
        RECT 105.480 38.270 105.620 44.070 ;
        RECT 107.320 43.370 107.460 47.050 ;
        RECT 107.260 43.050 107.520 43.370 ;
        RECT 109.620 41.670 109.760 66.510 ;
        RECT 111.000 64.110 111.140 68.550 ;
        RECT 115.080 67.870 115.340 68.190 ;
        RECT 115.140 66.830 115.280 67.870 ;
        RECT 115.080 66.510 115.340 66.830 ;
        RECT 113.230 64.275 114.770 64.645 ;
        RECT 110.940 63.790 111.200 64.110 ;
        RECT 111.000 58.670 111.140 63.790 ;
        RECT 112.780 62.770 113.040 63.090 ;
        RECT 110.940 58.350 111.200 58.670 ;
        RECT 110.480 54.270 110.740 54.590 ;
        RECT 110.020 51.890 110.280 52.210 ;
        RECT 110.080 47.790 110.220 51.890 ;
        RECT 110.540 50.510 110.680 54.270 ;
        RECT 112.840 52.550 112.980 62.770 ;
        RECT 113.700 62.430 113.960 62.750 ;
        RECT 114.160 62.430 114.420 62.750 ;
        RECT 113.760 60.710 113.900 62.430 ;
        RECT 114.220 61.390 114.360 62.430 ;
        RECT 114.160 61.070 114.420 61.390 ;
        RECT 115.600 61.050 115.740 74.670 ;
        RECT 118.360 74.310 118.500 76.710 ;
        RECT 118.820 74.990 118.960 82.490 ;
        RECT 121.520 81.130 121.780 81.450 ;
        RECT 119.220 79.090 119.480 79.410 ;
        RECT 118.760 74.670 119.020 74.990 ;
        RECT 119.280 74.650 119.420 79.090 ;
        RECT 121.060 78.410 121.320 78.730 ;
        RECT 121.120 77.030 121.260 78.410 ;
        RECT 121.580 77.710 121.720 81.130 ;
        RECT 122.040 77.710 122.180 82.490 ;
        RECT 122.440 81.130 122.700 81.450 ;
        RECT 122.500 79.070 122.640 81.130 ;
        RECT 122.960 80.430 123.100 83.850 ;
        RECT 124.800 82.130 124.940 83.850 ;
        RECT 125.720 82.810 125.860 84.870 ;
        RECT 126.120 84.530 126.380 84.850 ;
        RECT 125.660 82.490 125.920 82.810 ;
        RECT 124.740 81.810 125.000 82.130 ;
        RECT 122.900 80.110 123.160 80.430 ;
        RECT 125.720 80.390 125.860 82.490 ;
        RECT 124.340 80.250 125.860 80.390 ;
        RECT 124.340 79.410 124.480 80.250 ;
        RECT 124.280 79.090 124.540 79.410 ;
        RECT 122.440 78.750 122.700 79.070 ;
        RECT 121.520 77.390 121.780 77.710 ;
        RECT 121.980 77.390 122.240 77.710 ;
        RECT 121.060 76.710 121.320 77.030 ;
        RECT 121.120 76.430 121.260 76.710 ;
        RECT 121.120 76.290 122.180 76.430 ;
        RECT 121.520 75.690 121.780 76.010 ;
        RECT 119.220 74.330 119.480 74.650 ;
        RECT 118.300 73.990 118.560 74.310 ;
        RECT 116.530 72.435 118.070 72.805 ;
        RECT 118.360 71.250 118.500 73.990 ;
        RECT 118.760 72.970 119.020 73.290 ;
        RECT 118.820 71.930 118.960 72.970 ;
        RECT 118.760 71.610 119.020 71.930 ;
        RECT 118.300 70.930 118.560 71.250 ;
        RECT 118.360 69.550 118.500 70.930 ;
        RECT 119.280 70.910 119.420 74.330 ;
        RECT 121.580 73.970 121.720 75.690 ;
        RECT 122.040 73.970 122.180 76.290 ;
        RECT 120.600 73.650 120.860 73.970 ;
        RECT 121.520 73.650 121.780 73.970 ;
        RECT 121.980 73.650 122.240 73.970 ;
        RECT 122.440 73.650 122.700 73.970 ;
        RECT 120.660 71.590 120.800 73.650 ;
        RECT 120.600 71.270 120.860 71.590 ;
        RECT 119.220 70.590 119.480 70.910 ;
        RECT 118.300 69.230 118.560 69.550 ;
        RECT 120.660 68.270 120.800 71.270 ;
        RECT 122.500 71.250 122.640 73.650 ;
        RECT 122.440 70.930 122.700 71.250 ;
        RECT 122.500 68.530 122.640 70.930 ;
        RECT 120.660 68.130 121.260 68.270 ;
        RECT 122.440 68.210 122.700 68.530 ;
        RECT 121.120 67.850 121.260 68.130 ;
        RECT 121.060 67.530 121.320 67.850 ;
        RECT 116.530 66.995 118.070 67.365 ;
        RECT 121.120 63.430 121.260 67.530 ;
        RECT 122.500 66.830 122.640 68.210 ;
        RECT 122.440 66.510 122.700 66.830 ;
        RECT 124.340 66.150 124.480 79.090 ;
        RECT 126.180 79.070 126.320 84.530 ;
        RECT 127.500 83.850 127.760 84.170 ;
        RECT 127.560 80.090 127.700 83.850 ;
        RECT 131.825 83.315 133.365 83.685 ;
        RECT 127.960 82.490 128.220 82.810 ;
        RECT 128.020 80.430 128.160 82.490 ;
        RECT 133.940 82.150 134.200 82.470 ;
        RECT 128.525 80.595 130.065 80.965 ;
        RECT 134.000 80.430 134.140 82.150 ;
        RECT 136.240 81.810 136.500 82.130 ;
        RECT 134.860 81.470 135.120 81.790 ;
        RECT 127.960 80.110 128.220 80.430 ;
        RECT 133.940 80.110 134.200 80.430 ;
        RECT 127.500 79.770 127.760 80.090 ;
        RECT 134.920 79.410 135.060 81.470 ;
        RECT 136.300 79.410 136.440 81.810 ;
        RECT 137.160 81.130 137.420 81.450 ;
        RECT 126.120 78.750 126.380 79.070 ;
        RECT 127.490 78.895 127.770 79.265 ;
        RECT 131.180 79.090 131.440 79.410 ;
        RECT 134.860 79.320 135.120 79.410 ;
        RECT 134.460 79.180 135.120 79.320 ;
        RECT 127.500 78.750 127.760 78.895 ;
        RECT 130.720 78.750 130.980 79.070 ;
        RECT 127.560 76.690 127.700 78.750 ;
        RECT 127.500 76.370 127.760 76.690 ;
        RECT 127.040 75.690 127.300 76.010 ;
        RECT 127.100 73.630 127.240 75.690 ;
        RECT 128.525 75.155 130.065 75.525 ;
        RECT 130.780 74.990 130.920 78.750 ;
        RECT 131.240 76.690 131.380 79.090 ;
        RECT 133.710 78.585 133.970 78.730 ;
        RECT 133.710 78.410 134.210 78.585 ;
        RECT 133.770 78.330 134.210 78.410 ;
        RECT 131.825 77.875 133.365 78.245 ;
        RECT 133.930 78.215 134.210 78.330 ;
        RECT 134.460 77.790 134.600 79.180 ;
        RECT 134.860 79.090 135.120 79.180 ;
        RECT 136.240 79.320 136.500 79.410 ;
        RECT 136.240 79.180 136.900 79.320 ;
        RECT 136.240 79.090 136.500 79.180 ;
        RECT 135.320 78.410 135.580 78.730 ;
        RECT 133.020 77.620 133.280 77.710 ;
        RECT 133.540 77.650 134.600 77.790 ;
        RECT 133.540 77.620 133.680 77.650 ;
        RECT 133.020 77.480 133.680 77.620 ;
        RECT 133.020 77.390 133.280 77.480 ;
        RECT 135.380 77.030 135.520 78.410 ;
        RECT 136.230 78.215 136.510 78.585 ;
        RECT 135.780 77.390 136.040 77.710 ;
        RECT 133.480 76.710 133.740 77.030 ;
        RECT 135.320 76.710 135.580 77.030 ;
        RECT 131.180 76.370 131.440 76.690 ;
        RECT 130.720 74.670 130.980 74.990 ;
        RECT 133.540 73.630 133.680 76.710 ;
        RECT 135.840 74.650 135.980 77.390 ;
        RECT 136.300 77.030 136.440 78.215 ;
        RECT 136.760 77.710 136.900 79.180 ;
        RECT 137.220 78.730 137.360 81.130 ;
        RECT 137.620 80.110 137.880 80.430 ;
        RECT 140.440 80.390 140.580 87.590 ;
        RECT 145.900 86.910 146.160 87.230 ;
        RECT 143.820 86.035 145.360 86.405 ;
        RECT 143.600 84.530 143.860 84.850 ;
        RECT 143.660 83.150 143.800 84.530 ;
        RECT 145.440 83.850 145.700 84.170 ;
        RECT 143.600 82.830 143.860 83.150 ;
        RECT 142.680 82.150 142.940 82.470 ;
        RECT 142.740 80.390 142.880 82.150 ;
        RECT 143.820 80.595 145.360 80.965 ;
        RECT 145.500 80.430 145.640 83.850 ;
        RECT 145.960 82.470 146.100 86.910 ;
        RECT 147.120 83.315 148.660 83.685 ;
        RECT 145.900 82.150 146.160 82.470 ;
        RECT 139.980 80.250 140.580 80.390 ;
        RECT 140.900 80.250 142.880 80.390 ;
        RECT 137.160 78.410 137.420 78.730 ;
        RECT 136.700 77.390 136.960 77.710 ;
        RECT 137.680 77.620 137.820 80.110 ;
        RECT 137.220 77.480 137.820 77.620 ;
        RECT 136.240 76.710 136.500 77.030 ;
        RECT 137.220 74.900 137.360 77.480 ;
        RECT 137.620 76.710 137.880 77.030 ;
        RECT 136.760 74.760 137.360 74.900 ;
        RECT 135.780 74.330 136.040 74.650 ;
        RECT 127.040 73.310 127.300 73.630 ;
        RECT 127.500 73.310 127.760 73.630 ;
        RECT 133.480 73.310 133.740 73.630 ;
        RECT 127.100 71.590 127.240 73.310 ;
        RECT 127.560 71.930 127.700 73.310 ;
        RECT 131.825 72.435 133.365 72.805 ;
        RECT 127.500 71.610 127.760 71.930 ;
        RECT 127.040 71.270 127.300 71.590 ;
        RECT 124.280 65.830 124.540 66.150 ;
        RECT 122.440 64.810 122.700 65.130 ;
        RECT 122.500 64.110 122.640 64.810 ;
        RECT 122.440 63.790 122.700 64.110 ;
        RECT 121.060 63.110 121.320 63.430 ;
        RECT 116.530 61.555 118.070 61.925 ;
        RECT 115.540 60.730 115.800 61.050 ;
        RECT 113.700 60.390 113.960 60.710 ;
        RECT 113.230 58.835 114.770 59.205 ;
        RECT 120.600 57.330 120.860 57.650 ;
        RECT 118.300 56.650 118.560 56.970 ;
        RECT 116.530 56.115 118.070 56.485 ;
        RECT 118.360 55.270 118.500 56.650 ;
        RECT 115.080 54.950 115.340 55.270 ;
        RECT 118.300 54.950 118.560 55.270 ;
        RECT 113.230 53.395 114.770 53.765 ;
        RECT 110.940 52.230 111.200 52.550 ;
        RECT 112.780 52.230 113.040 52.550 ;
        RECT 110.480 50.190 110.740 50.510 ;
        RECT 110.020 47.470 110.280 47.790 ;
        RECT 110.540 45.070 110.680 50.190 ;
        RECT 111.000 48.810 111.140 52.230 ;
        RECT 111.400 51.890 111.660 52.210 ;
        RECT 110.940 48.490 111.200 48.810 ;
        RECT 111.000 47.790 111.140 48.490 ;
        RECT 111.460 47.790 111.600 51.890 ;
        RECT 115.140 51.870 115.280 54.950 ;
        RECT 115.540 53.930 115.800 54.250 ;
        RECT 118.300 53.930 118.560 54.250 ;
        RECT 120.140 53.930 120.400 54.250 ;
        RECT 115.600 53.230 115.740 53.930 ;
        RECT 118.360 53.230 118.500 53.930 ;
        RECT 115.540 52.910 115.800 53.230 ;
        RECT 118.300 52.910 118.560 53.230 ;
        RECT 120.200 52.210 120.340 53.930 ;
        RECT 120.140 51.890 120.400 52.210 ;
        RECT 112.320 51.550 112.580 51.870 ;
        RECT 115.080 51.550 115.340 51.870 ;
        RECT 111.860 49.170 112.120 49.490 ;
        RECT 110.940 47.470 111.200 47.790 ;
        RECT 111.400 47.470 111.660 47.790 ;
        RECT 111.920 45.070 112.060 49.170 ;
        RECT 112.380 45.830 112.520 51.550 ;
        RECT 116.530 50.675 118.070 51.045 ;
        RECT 115.080 49.850 115.340 50.170 ;
        RECT 113.230 47.955 114.770 48.325 ;
        RECT 112.380 45.690 113.440 45.830 ;
        RECT 110.480 44.750 110.740 45.070 ;
        RECT 111.860 44.750 112.120 45.070 ;
        RECT 109.560 41.350 109.820 41.670 ;
        RECT 106.340 39.310 106.600 39.630 ;
        RECT 105.420 37.950 105.680 38.270 ;
        RECT 104.960 37.610 105.220 37.930 ;
        RECT 105.020 34.190 105.160 37.610 ;
        RECT 104.960 33.870 105.220 34.190 ;
        RECT 102.660 33.450 103.780 33.510 ;
        RECT 102.660 33.190 102.920 33.450 ;
        RECT 104.040 33.190 104.300 33.510 ;
        RECT 102.200 32.170 102.460 32.490 ;
        RECT 105.020 32.230 105.160 33.870 ;
        RECT 105.480 32.830 105.620 37.950 ;
        RECT 105.880 35.910 106.140 36.230 ;
        RECT 105.940 34.190 106.080 35.910 ;
        RECT 106.400 34.190 106.540 39.310 ;
        RECT 107.260 38.630 107.520 38.950 ;
        RECT 109.560 38.630 109.820 38.950 ;
        RECT 110.020 38.630 110.280 38.950 ;
        RECT 107.320 35.890 107.460 38.630 ;
        RECT 109.620 36.910 109.760 38.630 ;
        RECT 109.560 36.590 109.820 36.910 ;
        RECT 107.260 35.570 107.520 35.890 ;
        RECT 109.560 35.570 109.820 35.890 ;
        RECT 105.880 33.870 106.140 34.190 ;
        RECT 106.340 33.870 106.600 34.190 ;
        RECT 105.880 33.190 106.140 33.510 ;
        RECT 105.940 32.830 106.080 33.190 ;
        RECT 107.720 32.850 107.980 33.170 ;
        RECT 105.420 32.510 105.680 32.830 ;
        RECT 105.880 32.510 106.140 32.830 ;
        RECT 105.940 32.230 106.080 32.510 ;
        RECT 105.020 32.090 106.080 32.230 ;
        RECT 107.780 31.470 107.920 32.850 ;
        RECT 109.620 32.830 109.760 35.570 ;
        RECT 110.080 34.190 110.220 38.630 ;
        RECT 111.920 38.270 112.060 44.750 ;
        RECT 113.300 44.730 113.440 45.690 ;
        RECT 115.140 45.070 115.280 49.850 ;
        RECT 120.140 47.470 120.400 47.790 ;
        RECT 116.530 45.235 118.070 45.605 ;
        RECT 115.080 44.750 115.340 45.070 ;
        RECT 113.240 44.410 113.500 44.730 ;
        RECT 120.200 44.390 120.340 47.470 ;
        RECT 120.660 46.090 120.800 57.330 ;
        RECT 120.600 45.770 120.860 46.090 ;
        RECT 120.140 44.070 120.400 44.390 ;
        RECT 113.230 42.515 114.770 42.885 ;
        RECT 116.530 39.795 118.070 40.165 ;
        RECT 121.120 39.540 121.260 63.110 ;
        RECT 121.980 62.090 122.240 62.410 ;
        RECT 126.120 62.090 126.380 62.410 ;
        RECT 122.040 61.390 122.180 62.090 ;
        RECT 121.980 61.070 122.240 61.390 ;
        RECT 123.820 59.370 124.080 59.690 ;
        RECT 123.880 57.650 124.020 59.370 ;
        RECT 126.180 57.650 126.320 62.090 ;
        RECT 127.100 60.710 127.240 71.270 ;
        RECT 133.540 70.570 133.680 73.310 ;
        RECT 135.320 72.970 135.580 73.290 ;
        RECT 134.400 71.270 134.660 71.590 ;
        RECT 127.500 70.250 127.760 70.570 ;
        RECT 133.480 70.250 133.740 70.570 ;
        RECT 127.560 65.810 127.700 70.250 ;
        RECT 128.525 69.715 130.065 70.085 ;
        RECT 134.460 69.550 134.600 71.270 ;
        RECT 135.380 69.550 135.520 72.970 ;
        RECT 136.760 72.270 136.900 74.760 ;
        RECT 137.680 73.970 137.820 76.710 ;
        RECT 139.000 75.690 139.260 76.010 ;
        RECT 139.060 74.990 139.200 75.690 ;
        RECT 139.000 74.670 139.260 74.990 ;
        RECT 138.080 73.990 138.340 74.310 ;
        RECT 137.620 73.650 137.880 73.970 ;
        RECT 136.700 71.950 136.960 72.270 ;
        RECT 137.620 71.270 137.880 71.590 ;
        RECT 134.400 69.230 134.660 69.550 ;
        RECT 135.320 69.230 135.580 69.550 ;
        RECT 131.825 66.995 133.365 67.365 ;
        RECT 127.960 66.170 128.220 66.490 ;
        RECT 127.500 65.490 127.760 65.810 ;
        RECT 128.020 64.110 128.160 66.170 ;
        RECT 134.460 66.150 134.600 69.230 ;
        RECT 137.680 69.210 137.820 71.270 ;
        RECT 138.140 69.550 138.280 73.990 ;
        RECT 139.060 72.270 139.200 74.670 ;
        RECT 139.000 71.950 139.260 72.270 ;
        RECT 138.540 70.590 138.800 70.910 ;
        RECT 138.600 69.550 138.740 70.590 ;
        RECT 138.080 69.230 138.340 69.550 ;
        RECT 138.540 69.230 138.800 69.550 ;
        RECT 137.620 68.890 137.880 69.210 ;
        RECT 135.320 67.530 135.580 67.850 ;
        RECT 134.400 65.830 134.660 66.150 ;
        RECT 135.380 65.810 135.520 67.530 ;
        RECT 138.140 66.830 138.280 69.230 ;
        RECT 138.080 66.510 138.340 66.830 ;
        RECT 139.980 66.150 140.120 80.250 ;
        RECT 140.900 79.265 141.040 80.250 ;
        RECT 145.440 80.110 145.700 80.430 ;
        RECT 140.830 78.895 141.110 79.265 ;
        RECT 143.140 78.410 143.400 78.730 ;
        RECT 140.380 76.710 140.640 77.030 ;
        RECT 140.440 72.270 140.580 76.710 ;
        RECT 143.200 76.690 143.340 78.410 ;
        RECT 145.500 77.710 145.640 80.110 ;
        RECT 145.960 79.410 146.100 82.150 ;
        RECT 145.900 79.090 146.160 79.410 ;
        RECT 145.440 77.390 145.700 77.710 ;
        RECT 143.140 76.370 143.400 76.690 ;
        RECT 141.300 75.690 141.560 76.010 ;
        RECT 141.760 75.690 142.020 76.010 ;
        RECT 142.680 75.690 142.940 76.010 ;
        RECT 141.360 74.990 141.500 75.690 ;
        RECT 141.300 74.670 141.560 74.990 ;
        RECT 141.300 73.650 141.560 73.970 ;
        RECT 140.840 72.970 141.100 73.290 ;
        RECT 140.380 71.950 140.640 72.270 ;
        RECT 140.440 71.250 140.580 71.950 ;
        RECT 140.380 70.930 140.640 71.250 ;
        RECT 140.900 70.910 141.040 72.970 ;
        RECT 140.840 70.590 141.100 70.910 ;
        RECT 140.380 70.250 140.640 70.570 ;
        RECT 140.440 69.550 140.580 70.250 ;
        RECT 140.380 69.230 140.640 69.550 ;
        RECT 140.840 68.550 141.100 68.870 ;
        RECT 139.920 65.830 140.180 66.150 ;
        RECT 135.320 65.490 135.580 65.810 ;
        RECT 140.900 65.130 141.040 68.550 ;
        RECT 141.360 65.470 141.500 73.650 ;
        RECT 141.820 68.530 141.960 75.690 ;
        RECT 142.740 74.650 142.880 75.690 ;
        RECT 142.680 74.330 142.940 74.650 ;
        RECT 143.200 73.970 143.340 76.370 ;
        RECT 145.440 75.690 145.700 76.010 ;
        RECT 143.820 75.155 145.360 75.525 ;
        RECT 142.220 73.650 142.480 73.970 ;
        RECT 143.140 73.650 143.400 73.970 ;
        RECT 143.600 73.650 143.860 73.970 ;
        RECT 141.760 68.210 142.020 68.530 ;
        RECT 142.280 65.810 142.420 73.650 ;
        RECT 143.140 72.970 143.400 73.290 ;
        RECT 143.200 71.590 143.340 72.970 ;
        RECT 143.140 71.270 143.400 71.590 ;
        RECT 143.660 71.250 143.800 73.650 ;
        RECT 145.500 72.270 145.640 75.690 ;
        RECT 145.960 73.970 146.100 79.090 ;
        RECT 147.120 77.875 148.660 78.245 ;
        RECT 146.820 75.690 147.080 76.010 ;
        RECT 146.880 74.990 147.020 75.690 ;
        RECT 146.820 74.670 147.080 74.990 ;
        RECT 145.900 73.650 146.160 73.970 ;
        RECT 146.360 73.650 146.620 73.970 ;
        RECT 145.900 72.970 146.160 73.290 ;
        RECT 145.440 71.950 145.700 72.270 ;
        RECT 142.680 70.930 142.940 71.250 ;
        RECT 143.600 70.930 143.860 71.250 ;
        RECT 145.500 70.990 145.640 71.950 ;
        RECT 145.960 71.590 146.100 72.970 ;
        RECT 145.900 71.270 146.160 71.590 ;
        RECT 142.740 67.850 142.880 70.930 ;
        RECT 143.140 70.590 143.400 70.910 ;
        RECT 145.500 70.850 146.100 70.990 ;
        RECT 143.200 68.950 143.340 70.590 ;
        RECT 145.440 70.250 145.700 70.570 ;
        RECT 143.820 69.715 145.360 70.085 ;
        RECT 144.060 69.230 144.320 69.550 ;
        RECT 143.200 68.870 143.800 68.950 ;
        RECT 143.200 68.810 143.860 68.870 ;
        RECT 143.600 68.550 143.860 68.810 ;
        RECT 143.140 68.210 143.400 68.530 ;
        RECT 142.680 67.530 142.940 67.850 ;
        RECT 143.200 66.830 143.340 68.210 ;
        RECT 143.140 66.510 143.400 66.830 ;
        RECT 144.120 66.150 144.260 69.230 ;
        RECT 145.500 68.870 145.640 70.250 ;
        RECT 145.440 68.550 145.700 68.870 ;
        RECT 145.960 68.270 146.100 70.850 ;
        RECT 146.420 69.550 146.560 73.650 ;
        RECT 147.120 72.435 148.660 72.805 ;
        RECT 148.660 71.610 148.920 71.930 ;
        RECT 146.820 71.270 147.080 71.590 ;
        RECT 147.280 71.270 147.540 71.590 ;
        RECT 146.360 69.230 146.620 69.550 ;
        RECT 146.880 68.950 147.020 71.270 ;
        RECT 145.040 68.130 146.100 68.270 ;
        RECT 146.420 68.810 147.020 68.950 ;
        RECT 145.040 67.850 145.180 68.130 ;
        RECT 144.980 67.530 145.240 67.850 ;
        RECT 145.440 67.530 145.700 67.850 ;
        RECT 145.900 67.530 146.160 67.850 ;
        RECT 145.500 66.150 145.640 67.530 ;
        RECT 145.960 66.150 146.100 67.530 ;
        RECT 144.060 65.830 144.320 66.150 ;
        RECT 145.440 65.830 145.700 66.150 ;
        RECT 145.900 65.830 146.160 66.150 ;
        RECT 142.220 65.490 142.480 65.810 ;
        RECT 141.300 65.150 141.560 65.470 ;
        RECT 142.740 65.410 144.260 65.550 ;
        RECT 142.740 65.130 142.880 65.410 ;
        RECT 144.120 65.130 144.260 65.410 ;
        RECT 138.080 64.810 138.340 65.130 ;
        RECT 140.840 64.810 141.100 65.130 ;
        RECT 142.680 64.810 142.940 65.130 ;
        RECT 143.140 64.810 143.400 65.130 ;
        RECT 144.060 64.810 144.320 65.130 ;
        RECT 128.525 64.275 130.065 64.645 ;
        RECT 127.960 63.790 128.220 64.110 ;
        RECT 131.825 61.555 133.365 61.925 ;
        RECT 138.140 61.390 138.280 64.810 ;
        RECT 143.200 63.770 143.340 64.810 ;
        RECT 143.820 64.275 145.360 64.645 ;
        RECT 143.140 63.450 143.400 63.770 ;
        RECT 142.680 62.090 142.940 62.410 ;
        RECT 138.080 61.070 138.340 61.390 ;
        RECT 127.040 60.390 127.300 60.710 ;
        RECT 123.820 57.330 124.080 57.650 ;
        RECT 126.120 57.330 126.380 57.650 ;
        RECT 125.660 56.650 125.920 56.970 ;
        RECT 125.720 55.610 125.860 56.650 ;
        RECT 125.660 55.290 125.920 55.610 ;
        RECT 121.980 53.930 122.240 54.250 ;
        RECT 122.040 52.210 122.180 53.930 ;
        RECT 121.980 51.890 122.240 52.210 ;
        RECT 121.520 51.550 121.780 51.870 ;
        RECT 121.580 50.510 121.720 51.550 ;
        RECT 121.520 50.190 121.780 50.510 ;
        RECT 122.040 50.170 122.180 51.890 ;
        RECT 122.440 51.210 122.700 51.530 ;
        RECT 121.980 49.850 122.240 50.170 ;
        RECT 122.040 39.630 122.180 49.850 ;
        RECT 121.520 39.540 121.780 39.630 ;
        RECT 121.120 39.400 121.780 39.540 ;
        RECT 121.520 39.310 121.780 39.400 ;
        RECT 121.980 39.310 122.240 39.630 ;
        RECT 115.540 38.970 115.800 39.290 ;
        RECT 122.500 39.030 122.640 51.210 ;
        RECT 126.180 46.510 126.320 57.330 ;
        RECT 126.180 46.430 126.780 46.510 ;
        RECT 126.180 46.370 126.840 46.430 ;
        RECT 126.580 46.110 126.840 46.370 ;
        RECT 127.100 44.730 127.240 60.390 ;
        RECT 128.525 58.835 130.065 59.205 ;
        RECT 142.740 57.990 142.880 62.090 ;
        RECT 143.820 58.835 145.360 59.205 ;
        RECT 131.180 57.670 131.440 57.990 ;
        RECT 142.680 57.670 142.940 57.990 ;
        RECT 127.960 57.330 128.220 57.650 ;
        RECT 127.500 56.650 127.760 56.970 ;
        RECT 127.560 55.950 127.700 56.650 ;
        RECT 127.500 55.630 127.760 55.950 ;
        RECT 128.020 53.230 128.160 57.330 ;
        RECT 130.260 56.990 130.520 57.310 ;
        RECT 128.525 53.395 130.065 53.765 ;
        RECT 127.960 52.910 128.220 53.230 ;
        RECT 130.320 52.210 130.460 56.990 ;
        RECT 130.720 54.950 130.980 55.270 ;
        RECT 130.780 52.210 130.920 54.950 ;
        RECT 131.240 52.210 131.380 57.670 ;
        RECT 135.320 57.330 135.580 57.650 ;
        RECT 141.300 57.330 141.560 57.650 ;
        RECT 133.480 56.650 133.740 56.970 ;
        RECT 131.825 56.115 133.365 56.485 ;
        RECT 133.540 55.610 133.680 56.650 ;
        RECT 133.480 55.290 133.740 55.610 ;
        RECT 133.480 52.910 133.740 53.230 ;
        RECT 130.260 51.890 130.520 52.210 ;
        RECT 130.720 51.890 130.980 52.210 ;
        RECT 131.180 51.890 131.440 52.210 ;
        RECT 127.500 51.210 127.760 51.530 ;
        RECT 127.560 50.510 127.700 51.210 ;
        RECT 127.500 50.190 127.760 50.510 ;
        RECT 128.880 50.190 129.140 50.510 ;
        RECT 128.940 49.490 129.080 50.190 ;
        RECT 128.880 49.170 129.140 49.490 ;
        RECT 128.525 47.955 130.065 48.325 ;
        RECT 129.340 47.130 129.600 47.450 ;
        RECT 129.400 45.070 129.540 47.130 ;
        RECT 130.780 47.110 130.920 51.890 ;
        RECT 131.825 50.675 133.365 51.045 ;
        RECT 131.180 49.850 131.440 50.170 ;
        RECT 130.720 46.790 130.980 47.110 ;
        RECT 131.240 45.070 131.380 49.850 ;
        RECT 133.540 49.830 133.680 52.910 ;
        RECT 135.380 52.550 135.520 57.330 ;
        RECT 136.240 56.990 136.500 57.310 ;
        RECT 136.300 54.250 136.440 56.990 ;
        RECT 141.360 55.610 141.500 57.330 ;
        RECT 141.300 55.290 141.560 55.610 ;
        RECT 136.240 53.930 136.500 54.250 ;
        RECT 135.320 52.230 135.580 52.550 ;
        RECT 134.400 51.950 134.660 52.210 ;
        RECT 134.000 51.890 134.660 51.950 ;
        RECT 134.860 51.890 135.120 52.210 ;
        RECT 134.000 51.810 134.600 51.890 ;
        RECT 134.000 50.510 134.140 51.810 ;
        RECT 134.400 51.210 134.660 51.530 ;
        RECT 134.460 50.510 134.600 51.210 ;
        RECT 133.940 50.190 134.200 50.510 ;
        RECT 134.400 50.190 134.660 50.510 ;
        RECT 134.920 50.170 135.060 51.890 ;
        RECT 136.300 51.870 136.440 53.930 ;
        RECT 140.380 52.910 140.640 53.230 ;
        RECT 137.620 52.230 137.880 52.550 ;
        RECT 136.240 51.780 136.500 51.870 ;
        RECT 135.840 51.640 136.500 51.780 ;
        RECT 135.840 50.510 135.980 51.640 ;
        RECT 136.240 51.550 136.500 51.640 ;
        RECT 135.780 50.190 136.040 50.510 ;
        RECT 137.680 50.170 137.820 52.230 ;
        RECT 138.540 51.210 138.800 51.530 ;
        RECT 138.600 50.510 138.740 51.210 ;
        RECT 138.540 50.190 138.800 50.510 ;
        RECT 134.860 49.850 135.120 50.170 ;
        RECT 137.620 49.850 137.880 50.170 ;
        RECT 133.480 49.510 133.740 49.830 ;
        RECT 134.400 49.170 134.660 49.490 ;
        RECT 131.825 45.235 133.365 45.605 ;
        RECT 134.460 45.070 134.600 49.170 ;
        RECT 134.920 45.070 135.060 49.850 ;
        RECT 129.340 44.750 129.600 45.070 ;
        RECT 131.180 44.750 131.440 45.070 ;
        RECT 134.400 44.750 134.660 45.070 ;
        RECT 134.860 44.750 135.120 45.070 ;
        RECT 127.040 44.410 127.300 44.730 ;
        RECT 139.000 44.410 139.260 44.730 ;
        RECT 140.440 44.470 140.580 52.910 ;
        RECT 141.360 52.210 141.500 55.290 ;
        RECT 142.680 54.610 142.940 54.930 ;
        RECT 141.300 51.890 141.560 52.210 ;
        RECT 140.840 44.470 141.100 44.730 ;
        RECT 140.440 44.410 141.100 44.470 ;
        RECT 127.960 44.070 128.220 44.390 ;
        RECT 131.640 44.070 131.900 44.390 ;
        RECT 127.040 43.730 127.300 44.050 ;
        RECT 126.580 43.050 126.840 43.370 ;
        RECT 112.320 38.290 112.580 38.610 ;
        RECT 111.860 37.950 112.120 38.270 ;
        RECT 110.940 37.610 111.200 37.930 ;
        RECT 111.400 37.610 111.660 37.930 ;
        RECT 111.000 36.910 111.140 37.610 ;
        RECT 110.940 36.590 111.200 36.910 ;
        RECT 110.940 35.570 111.200 35.890 ;
        RECT 110.020 33.870 110.280 34.190 ;
        RECT 109.560 32.510 109.820 32.830 ;
        RECT 111.000 32.490 111.140 35.570 ;
        RECT 111.460 34.190 111.600 37.610 ;
        RECT 111.920 35.890 112.060 37.950 ;
        RECT 111.860 35.570 112.120 35.890 ;
        RECT 111.400 33.870 111.660 34.190 ;
        RECT 111.400 33.420 111.660 33.510 ;
        RECT 111.920 33.420 112.060 35.570 ;
        RECT 112.380 33.510 112.520 38.290 ;
        RECT 112.770 38.095 113.050 38.465 ;
        RECT 115.080 38.290 115.340 38.610 ;
        RECT 112.780 37.950 113.040 38.095 ;
        RECT 113.230 37.075 114.770 37.445 ;
        RECT 112.780 35.910 113.040 36.230 ;
        RECT 112.840 33.510 112.980 35.910 ;
        RECT 114.620 34.890 114.880 35.210 ;
        RECT 114.680 33.510 114.820 34.890 ;
        RECT 115.140 34.190 115.280 38.290 ;
        RECT 115.600 36.230 115.740 38.970 ;
        RECT 119.280 38.950 122.640 39.030 ;
        RECT 119.280 38.890 122.700 38.950 ;
        RECT 116.000 38.290 116.260 38.610 ;
        RECT 117.840 38.290 118.100 38.610 ;
        RECT 116.060 36.570 116.200 38.290 ;
        RECT 117.900 37.785 118.040 38.290 ;
        RECT 117.830 37.415 118.110 37.785 ;
        RECT 118.760 37.610 119.020 37.930 ;
        RECT 116.000 36.250 116.260 36.570 ;
        RECT 115.540 35.910 115.800 36.230 ;
        RECT 115.080 33.870 115.340 34.190 ;
        RECT 115.600 33.510 115.740 35.910 ;
        RECT 116.000 35.570 116.260 35.890 ;
        RECT 116.060 33.850 116.200 35.570 ;
        RECT 116.530 34.355 118.070 34.725 ;
        RECT 118.820 34.190 118.960 37.610 ;
        RECT 119.280 35.890 119.420 38.890 ;
        RECT 119.680 38.290 119.940 38.610 ;
        RECT 119.740 36.910 119.880 38.290 ;
        RECT 121.060 37.950 121.320 38.270 ;
        RECT 121.520 37.950 121.780 38.270 ;
        RECT 120.140 37.610 120.400 37.930 ;
        RECT 119.680 36.590 119.940 36.910 ;
        RECT 120.200 36.570 120.340 37.610 ;
        RECT 121.120 36.910 121.260 37.950 ;
        RECT 121.060 36.590 121.320 36.910 ;
        RECT 120.140 36.250 120.400 36.570 ;
        RECT 121.580 36.310 121.720 37.950 ;
        RECT 121.120 36.230 121.720 36.310 ;
        RECT 122.040 36.230 122.180 38.890 ;
        RECT 122.440 38.630 122.700 38.890 ;
        RECT 123.360 38.630 123.620 38.950 ;
        RECT 124.280 38.630 124.540 38.950 ;
        RECT 125.660 38.630 125.920 38.950 ;
        RECT 126.120 38.630 126.380 38.950 ;
        RECT 123.420 37.930 123.560 38.630 ;
        RECT 123.360 37.610 123.620 37.930 ;
        RECT 124.340 36.230 124.480 38.630 ;
        RECT 125.720 36.910 125.860 38.630 ;
        RECT 125.660 36.590 125.920 36.910 ;
        RECT 121.060 36.170 121.720 36.230 ;
        RECT 121.060 35.910 121.320 36.170 ;
        RECT 121.980 35.910 122.240 36.230 ;
        RECT 124.280 35.910 124.540 36.230 ;
        RECT 119.220 35.570 119.480 35.890 ;
        RECT 121.520 35.745 121.780 35.890 ;
        RECT 120.140 35.230 120.400 35.550 ;
        RECT 121.510 35.375 121.790 35.745 ;
        RECT 120.200 34.190 120.340 35.230 ;
        RECT 122.900 34.890 123.160 35.210 ;
        RECT 118.760 33.870 119.020 34.190 ;
        RECT 120.140 33.870 120.400 34.190 ;
        RECT 116.000 33.530 116.260 33.850 ;
        RECT 111.400 33.280 112.060 33.420 ;
        RECT 111.400 33.190 111.660 33.280 ;
        RECT 112.320 33.190 112.580 33.510 ;
        RECT 112.780 33.190 113.040 33.510 ;
        RECT 114.620 33.190 114.880 33.510 ;
        RECT 115.540 33.190 115.800 33.510 ;
        RECT 110.940 32.170 111.200 32.490 ;
        RECT 111.400 32.170 111.660 32.490 ;
        RECT 111.460 31.470 111.600 32.170 ;
        RECT 113.230 31.635 114.770 32.005 ;
        RECT 115.600 31.470 115.740 33.190 ;
        RECT 93.460 31.150 93.720 31.470 ;
        RECT 99.900 31.150 100.160 31.470 ;
        RECT 107.720 31.150 107.980 31.470 ;
        RECT 111.400 31.150 111.660 31.470 ;
        RECT 115.540 31.150 115.800 31.470 ;
        RECT 42.625 30.170 43.490 30.790 ;
        RECT 116.060 30.450 116.200 33.530 ;
        RECT 122.960 33.510 123.100 34.890 ;
        RECT 124.340 34.190 124.480 35.910 ;
        RECT 126.180 34.190 126.320 38.630 ;
        RECT 126.640 35.890 126.780 43.050 ;
        RECT 127.100 37.785 127.240 43.730 ;
        RECT 127.500 38.630 127.760 38.950 ;
        RECT 127.560 37.930 127.700 38.630 ;
        RECT 128.020 37.930 128.160 44.070 ;
        RECT 128.525 42.515 130.065 42.885 ;
        RECT 131.700 42.350 131.840 44.070 ;
        RECT 134.860 43.730 135.120 44.050 ;
        RECT 134.400 43.050 134.660 43.370 ;
        RECT 131.640 42.030 131.900 42.350 ;
        RECT 131.825 39.795 133.365 40.165 ;
        RECT 134.460 38.950 134.600 43.050 ;
        RECT 134.920 38.950 135.060 43.730 ;
        RECT 139.060 41.330 139.200 44.410 ;
        RECT 140.440 44.330 141.040 44.410 ;
        RECT 140.440 43.790 140.580 44.330 ;
        RECT 139.980 43.650 140.580 43.790 ;
        RECT 139.000 41.010 139.260 41.330 ;
        RECT 139.980 39.630 140.120 43.650 ;
        RECT 141.360 41.330 141.500 51.890 ;
        RECT 142.740 44.050 142.880 54.610 ;
        RECT 143.820 53.395 145.360 53.765 ;
        RECT 145.500 49.830 145.640 65.830 ;
        RECT 146.420 64.110 146.560 68.810 ;
        RECT 147.340 67.850 147.480 71.270 ;
        RECT 148.720 68.530 148.860 71.610 ;
        RECT 150.500 70.930 150.760 71.250 ;
        RECT 150.560 69.065 150.700 70.930 ;
        RECT 150.490 68.695 150.770 69.065 ;
        RECT 148.660 68.210 148.920 68.530 ;
        RECT 147.280 67.530 147.540 67.850 ;
        RECT 147.120 66.995 148.660 67.365 ;
        RECT 150.960 64.810 151.220 65.130 ;
        RECT 146.360 63.790 146.620 64.110 ;
        RECT 146.360 62.770 146.620 63.090 ;
        RECT 146.420 61.390 146.560 62.770 ;
        RECT 147.120 61.555 148.660 61.925 ;
        RECT 146.360 61.070 146.620 61.390 ;
        RECT 145.900 60.390 146.160 60.710 ;
        RECT 145.960 55.270 146.100 60.390 ;
        RECT 150.040 60.050 150.300 60.370 ;
        RECT 147.740 59.370 148.000 59.690 ;
        RECT 147.800 57.310 147.940 59.370 ;
        RECT 150.100 58.670 150.240 60.050 ;
        RECT 150.040 58.350 150.300 58.670 ;
        RECT 147.740 56.990 148.000 57.310 ;
        RECT 147.120 56.115 148.660 56.485 ;
        RECT 145.900 54.950 146.160 55.270 ;
        RECT 147.740 53.930 148.000 54.250 ;
        RECT 147.800 51.870 147.940 53.930 ;
        RECT 147.740 51.550 148.000 51.870 ;
        RECT 147.120 50.675 148.660 51.045 ;
        RECT 145.440 49.510 145.700 49.830 ;
        RECT 150.500 49.170 150.760 49.490 ;
        RECT 150.560 48.665 150.700 49.170 ;
        RECT 143.820 47.955 145.360 48.325 ;
        RECT 150.490 48.295 150.770 48.665 ;
        RECT 147.120 45.235 148.660 45.605 ;
        RECT 142.680 43.730 142.940 44.050 ;
        RECT 141.760 43.050 142.020 43.370 ;
        RECT 141.300 41.010 141.560 41.330 ;
        RECT 140.380 40.670 140.640 40.990 ;
        RECT 140.440 39.630 140.580 40.670 ;
        RECT 140.840 40.330 141.100 40.650 ;
        RECT 139.920 39.310 140.180 39.630 ;
        RECT 140.380 39.310 140.640 39.630 ;
        RECT 134.400 38.630 134.660 38.950 ;
        RECT 134.860 38.630 135.120 38.950 ;
        RECT 139.920 38.630 140.180 38.950 ;
        RECT 131.180 37.950 131.440 38.270 ;
        RECT 131.640 37.950 131.900 38.270 ;
        RECT 127.030 37.415 127.310 37.785 ;
        RECT 127.500 37.610 127.760 37.930 ;
        RECT 127.960 37.610 128.220 37.930 ;
        RECT 130.260 37.610 130.520 37.930 ;
        RECT 130.720 37.610 130.980 37.930 ;
        RECT 127.560 36.820 127.700 37.610 ;
        RECT 128.525 37.075 130.065 37.445 ;
        RECT 127.560 36.680 130.000 36.820 ;
        RECT 129.860 36.230 130.000 36.680 ;
        RECT 127.960 35.910 128.220 36.230 ;
        RECT 129.800 35.910 130.060 36.230 ;
        RECT 126.580 35.570 126.840 35.890 ;
        RECT 127.030 35.630 127.310 35.745 ;
        RECT 127.500 35.630 127.760 35.890 ;
        RECT 127.030 35.570 127.760 35.630 ;
        RECT 127.030 35.490 127.700 35.570 ;
        RECT 127.030 35.375 127.310 35.490 ;
        RECT 126.580 34.890 126.840 35.210 ;
        RECT 127.040 34.890 127.300 35.210 ;
        RECT 126.640 34.190 126.780 34.890 ;
        RECT 124.280 33.870 124.540 34.190 ;
        RECT 126.120 33.870 126.380 34.190 ;
        RECT 126.580 33.870 126.840 34.190 ;
        RECT 127.100 33.510 127.240 34.890 ;
        RECT 117.840 33.190 118.100 33.510 ;
        RECT 122.900 33.190 123.160 33.510 ;
        RECT 127.040 33.190 127.300 33.510 ;
        RECT 117.900 31.470 118.040 33.190 ;
        RECT 127.560 32.830 127.700 35.490 ;
        RECT 128.020 33.510 128.160 35.910 ;
        RECT 128.420 35.570 128.680 35.890 ;
        RECT 128.880 35.570 129.140 35.890 ;
        RECT 128.480 34.190 128.620 35.570 ;
        RECT 128.420 33.870 128.680 34.190 ;
        RECT 127.960 33.420 128.220 33.510 ;
        RECT 128.940 33.420 129.080 35.570 ;
        RECT 130.320 35.550 130.460 37.610 ;
        RECT 130.780 35.890 130.920 37.610 ;
        RECT 130.720 35.570 130.980 35.890 ;
        RECT 130.260 35.230 130.520 35.550 ;
        RECT 130.720 34.890 130.980 35.210 ;
        RECT 130.780 33.590 130.920 34.890 ;
        RECT 131.240 34.190 131.380 37.950 ;
        RECT 131.700 36.910 131.840 37.950 ;
        RECT 131.640 36.590 131.900 36.910 ;
        RECT 134.460 36.570 134.600 38.630 ;
        RECT 139.000 38.290 139.260 38.610 ;
        RECT 137.620 37.950 137.880 38.270 ;
        RECT 132.560 36.250 132.820 36.570 ;
        RECT 133.480 36.250 133.740 36.570 ;
        RECT 134.400 36.250 134.660 36.570 ;
        RECT 132.100 35.570 132.360 35.890 ;
        RECT 132.160 35.210 132.300 35.570 ;
        RECT 132.620 35.210 132.760 36.250 ;
        RECT 133.540 35.890 133.680 36.250 ;
        RECT 134.460 35.890 134.600 36.250 ;
        RECT 133.480 35.570 133.740 35.890 ;
        RECT 133.940 35.570 134.200 35.890 ;
        RECT 134.400 35.570 134.660 35.890 ;
        RECT 132.100 34.890 132.360 35.210 ;
        RECT 132.560 34.890 132.820 35.210 ;
        RECT 131.825 34.355 133.365 34.725 ;
        RECT 134.000 34.190 134.140 35.570 ;
        RECT 131.180 33.870 131.440 34.190 ;
        RECT 133.940 33.870 134.200 34.190 ;
        RECT 132.100 33.590 132.360 33.850 ;
        RECT 130.780 33.530 132.360 33.590 ;
        RECT 127.960 33.280 129.080 33.420 ;
        RECT 127.960 33.190 128.220 33.280 ;
        RECT 130.260 33.190 130.520 33.510 ;
        RECT 130.780 33.450 132.300 33.530 ;
        RECT 134.460 33.510 134.600 35.570 ;
        RECT 137.680 33.850 137.820 37.950 ;
        RECT 139.060 36.910 139.200 38.290 ;
        RECT 139.460 37.610 139.720 37.930 ;
        RECT 139.000 36.590 139.260 36.910 ;
        RECT 139.520 36.310 139.660 37.610 ;
        RECT 139.980 36.910 140.120 38.630 ;
        RECT 139.920 36.590 140.180 36.910 ;
        RECT 139.520 36.170 140.120 36.310 ;
        RECT 139.980 35.890 140.120 36.170 ;
        RECT 140.440 35.890 140.580 39.310 ;
        RECT 140.900 39.290 141.040 40.330 ;
        RECT 140.840 38.970 141.100 39.290 ;
        RECT 141.360 36.230 141.500 41.010 ;
        RECT 141.820 38.610 141.960 43.050 ;
        RECT 142.740 42.350 142.880 43.730 ;
        RECT 143.140 43.050 143.400 43.370 ;
        RECT 146.360 43.050 146.620 43.370 ;
        RECT 142.680 42.030 142.940 42.350 ;
        RECT 143.200 41.670 143.340 43.050 ;
        RECT 143.820 42.515 145.360 42.885 ;
        RECT 143.140 41.350 143.400 41.670 ;
        RECT 146.420 40.990 146.560 43.050 ;
        RECT 149.580 42.030 149.840 42.350 ;
        RECT 146.360 40.670 146.620 40.990 ;
        RECT 142.220 40.330 142.480 40.650 ;
        RECT 142.280 39.630 142.420 40.330 ;
        RECT 147.120 39.795 148.660 40.165 ;
        RECT 142.220 39.310 142.480 39.630 ;
        RECT 141.760 38.290 142.020 38.610 ;
        RECT 145.900 37.610 146.160 37.930 ;
        RECT 143.820 37.075 145.360 37.445 ;
        RECT 141.300 35.910 141.560 36.230 ;
        RECT 139.920 35.570 140.180 35.890 ;
        RECT 140.380 35.570 140.640 35.890 ;
        RECT 137.620 33.530 137.880 33.850 ;
        RECT 134.400 33.190 134.660 33.510 ;
        RECT 127.500 32.510 127.760 32.830 ;
        RECT 128.525 31.635 130.065 32.005 ;
        RECT 130.320 31.470 130.460 33.190 ;
        RECT 139.980 33.170 140.120 35.570 ;
        RECT 140.840 34.890 141.100 35.210 ;
        RECT 137.620 32.850 137.880 33.170 ;
        RECT 139.920 32.850 140.180 33.170 ;
        RECT 137.680 31.470 137.820 32.850 ;
        RECT 140.900 32.830 141.040 34.890 ;
        RECT 145.960 33.510 146.100 37.610 ;
        RECT 149.120 35.230 149.380 35.550 ;
        RECT 146.360 34.890 146.620 35.210 ;
        RECT 146.420 34.190 146.560 34.890 ;
        RECT 147.120 34.355 148.660 34.725 ;
        RECT 149.180 34.190 149.320 35.230 ;
        RECT 149.640 34.190 149.780 42.030 ;
        RECT 150.040 38.630 150.300 38.950 ;
        RECT 150.100 36.910 150.240 38.630 ;
        RECT 150.040 36.590 150.300 36.910 ;
        RECT 146.360 33.870 146.620 34.190 ;
        RECT 149.120 33.870 149.380 34.190 ;
        RECT 149.580 33.870 149.840 34.190 ;
        RECT 145.900 33.190 146.160 33.510 ;
        RECT 140.840 32.510 141.100 32.830 ;
        RECT 117.840 31.150 118.100 31.470 ;
        RECT 130.260 31.150 130.520 31.470 ;
        RECT 137.620 31.150 137.880 31.470 ;
        RECT 140.900 30.790 141.040 32.510 ;
        RECT 143.820 31.635 145.360 32.005 ;
        RECT 151.020 31.470 151.160 64.810 ;
        RECT 152.800 33.190 153.060 33.510 ;
        RECT 150.960 31.150 151.220 31.470 ;
        RECT 140.840 30.470 141.100 30.790 ;
        RECT 90.240 30.130 90.500 30.450 ;
        RECT 98.520 30.360 98.780 30.450 ;
        RECT 106.340 30.360 106.600 30.450 ;
        RECT 114.160 30.360 114.420 30.450 ;
        RECT 98.120 30.220 98.780 30.360 ;
        RECT 7.855 28.890 29.665 29.580 ;
        RECT 7.855 28.675 8.595 28.890 ;
        RECT 1.000 23.170 2.510 25.490 ;
        RECT 90.300 22.220 90.440 30.130 ;
        RECT 98.120 22.220 98.260 30.220 ;
        RECT 98.520 30.130 98.780 30.220 ;
        RECT 105.940 30.220 106.600 30.360 ;
        RECT 101.235 28.915 102.775 29.285 ;
        RECT 105.940 22.220 106.080 30.220 ;
        RECT 106.340 30.130 106.600 30.220 ;
        RECT 113.760 30.220 114.420 30.360 ;
        RECT 113.760 22.220 113.900 30.220 ;
        RECT 114.160 30.130 114.420 30.220 ;
        RECT 116.000 30.130 116.260 30.450 ;
        RECT 121.520 30.130 121.780 30.450 ;
        RECT 129.340 30.130 129.600 30.450 ;
        RECT 137.160 30.130 137.420 30.450 ;
        RECT 116.530 28.915 118.070 29.285 ;
        RECT 121.580 22.220 121.720 30.130 ;
        RECT 129.400 22.220 129.540 30.130 ;
        RECT 131.825 28.915 133.365 29.285 ;
        RECT 137.220 22.220 137.360 30.130 ;
        RECT 144.980 29.790 145.240 30.110 ;
        RECT 151.880 29.790 152.140 30.110 ;
        RECT 145.040 22.220 145.180 29.790 ;
        RECT 147.120 28.915 148.660 29.285 ;
        RECT 151.940 28.265 152.080 29.790 ;
        RECT 151.870 27.895 152.150 28.265 ;
        RECT 152.860 22.220 153.000 33.190 ;
        RECT 59.010 20.540 59.440 20.940 ;
        RECT 8.230 15.990 10.045 18.735 ;
        RECT 71.150 15.655 71.955 16.015 ;
        RECT 90.230 15.655 90.510 22.220 ;
        RECT 71.150 15.375 90.510 15.655 ;
        RECT 71.150 15.215 71.955 15.375 ;
        RECT 69.770 14.950 70.290 15.045 ;
        RECT 98.050 14.950 98.330 22.220 ;
        RECT 69.770 14.670 98.330 14.950 ;
        RECT 69.770 14.560 70.290 14.670 ;
        RECT 68.575 14.040 69.095 14.150 ;
        RECT 105.870 14.040 106.150 22.220 ;
        RECT 68.575 13.760 106.150 14.040 ;
        RECT 68.575 13.665 69.095 13.760 ;
        RECT 67.610 13.380 68.130 13.480 ;
        RECT 113.690 13.380 113.970 22.220 ;
        RECT 67.610 13.100 113.970 13.380 ;
        RECT 67.610 12.995 68.130 13.100 ;
        RECT 66.655 12.790 67.175 12.885 ;
        RECT 121.510 12.790 121.790 22.220 ;
        RECT 66.655 12.510 121.790 12.790 ;
        RECT 66.655 12.400 67.175 12.510 ;
        RECT 65.625 11.990 66.145 12.100 ;
        RECT 129.330 11.990 129.610 22.220 ;
        RECT 65.625 11.710 129.610 11.990 ;
        RECT 65.625 11.615 66.145 11.710 ;
        RECT 64.650 11.245 65.170 11.335 ;
        RECT 137.150 11.245 137.430 22.220 ;
        RECT 64.650 10.965 137.430 11.245 ;
        RECT 64.650 10.850 65.170 10.965 ;
        RECT 63.640 10.170 64.160 10.270 ;
        RECT 144.970 10.170 145.250 22.220 ;
        RECT 63.640 9.890 145.250 10.170 ;
        RECT 63.640 9.785 64.160 9.890 ;
        RECT 62.440 9.400 62.960 9.500 ;
        RECT 152.790 9.400 153.070 22.220 ;
        RECT 62.440 9.120 153.070 9.400 ;
        RECT 62.440 9.015 62.960 9.120 ;
        RECT 53.125 7.780 54.035 8.675 ;
        RECT 82.960 8.140 83.920 8.410 ;
        RECT 61.960 7.835 83.920 8.140 ;
        RECT 23.925 7.040 24.830 7.480 ;
        RECT 61.960 7.040 62.265 7.835 ;
        RECT 82.960 7.520 83.920 7.835 ;
        RECT 23.925 6.740 62.265 7.040 ;
        RECT 23.955 6.735 62.265 6.740 ;
      LAYER via2 ;
        RECT 84.935 222.570 85.235 222.870 ;
        RECT 88.605 222.575 88.905 222.875 ;
        RECT 5.140 211.425 5.455 211.705 ;
        RECT 147.350 220.825 147.950 221.425 ;
        RECT 157.250 220.850 157.800 221.400 ;
        RECT 143.660 218.960 144.260 219.560 ;
        RECT 156.005 218.985 156.555 219.535 ;
        RECT 139.980 216.780 140.580 217.380 ;
        RECT 153.650 216.805 154.200 217.355 ;
        RECT 136.320 215.115 136.920 215.715 ;
        RECT 153.890 215.140 154.440 215.690 ;
        RECT 3.615 207.490 3.910 207.775 ;
        RECT 1.495 194.185 1.995 194.685 ;
        RECT 76.545 194.290 76.825 194.570 ;
        RECT 76.945 194.290 77.225 194.570 ;
        RECT 77.345 194.290 77.625 194.570 ;
        RECT 77.745 194.290 78.025 194.570 ;
        RECT 88.620 194.290 88.900 194.570 ;
        RECT 89.020 194.290 89.300 194.570 ;
        RECT 89.420 194.290 89.700 194.570 ;
        RECT 89.820 194.290 90.100 194.570 ;
        RECT 100.695 194.290 100.975 194.570 ;
        RECT 101.095 194.290 101.375 194.570 ;
        RECT 101.495 194.290 101.775 194.570 ;
        RECT 101.895 194.290 102.175 194.570 ;
        RECT 112.770 194.290 113.050 194.570 ;
        RECT 113.170 194.290 113.450 194.570 ;
        RECT 113.570 194.290 113.850 194.570 ;
        RECT 113.970 194.290 114.250 194.570 ;
        RECT 79.845 191.570 80.125 191.850 ;
        RECT 80.245 191.570 80.525 191.850 ;
        RECT 80.645 191.570 80.925 191.850 ;
        RECT 81.045 191.570 81.325 191.850 ;
        RECT 70.420 189.190 70.700 189.470 ;
        RECT 76.545 188.850 76.825 189.130 ;
        RECT 76.945 188.850 77.225 189.130 ;
        RECT 77.345 188.850 77.625 189.130 ;
        RECT 77.745 188.850 78.025 189.130 ;
        RECT 91.920 191.570 92.200 191.850 ;
        RECT 92.320 191.570 92.600 191.850 ;
        RECT 92.720 191.570 93.000 191.850 ;
        RECT 93.120 191.570 93.400 191.850 ;
        RECT 79.845 186.130 80.125 186.410 ;
        RECT 80.245 186.130 80.525 186.410 ;
        RECT 80.645 186.130 80.925 186.410 ;
        RECT 81.045 186.130 81.325 186.410 ;
        RECT 76.545 183.410 76.825 183.690 ;
        RECT 76.945 183.410 77.225 183.690 ;
        RECT 77.345 183.410 77.625 183.690 ;
        RECT 77.745 183.410 78.025 183.690 ;
        RECT 76.545 177.970 76.825 178.250 ;
        RECT 76.945 177.970 77.225 178.250 ;
        RECT 77.345 177.970 77.625 178.250 ;
        RECT 77.745 177.970 78.025 178.250 ;
        RECT 79.845 180.690 80.125 180.970 ;
        RECT 80.245 180.690 80.525 180.970 ;
        RECT 80.645 180.690 80.925 180.970 ;
        RECT 81.045 180.690 81.325 180.970 ;
        RECT 79.845 175.250 80.125 175.530 ;
        RECT 80.245 175.250 80.525 175.530 ;
        RECT 80.645 175.250 80.925 175.530 ;
        RECT 81.045 175.250 81.325 175.530 ;
        RECT 76.545 172.530 76.825 172.810 ;
        RECT 76.945 172.530 77.225 172.810 ;
        RECT 77.345 172.530 77.625 172.810 ;
        RECT 77.745 172.530 78.025 172.810 ;
        RECT 79.845 169.810 80.125 170.090 ;
        RECT 80.245 169.810 80.525 170.090 ;
        RECT 80.645 169.810 80.925 170.090 ;
        RECT 81.045 169.810 81.325 170.090 ;
        RECT 76.545 167.090 76.825 167.370 ;
        RECT 76.945 167.090 77.225 167.370 ;
        RECT 77.345 167.090 77.625 167.370 ;
        RECT 77.745 167.090 78.025 167.370 ;
        RECT 79.845 164.370 80.125 164.650 ;
        RECT 80.245 164.370 80.525 164.650 ;
        RECT 80.645 164.370 80.925 164.650 ;
        RECT 81.045 164.370 81.325 164.650 ;
        RECT 76.545 161.650 76.825 161.930 ;
        RECT 76.945 161.650 77.225 161.930 ;
        RECT 77.345 161.650 77.625 161.930 ;
        RECT 77.745 161.650 78.025 161.930 ;
        RECT 79.845 158.930 80.125 159.210 ;
        RECT 80.245 158.930 80.525 159.210 ;
        RECT 80.645 158.930 80.925 159.210 ;
        RECT 81.045 158.930 81.325 159.210 ;
        RECT 76.545 156.210 76.825 156.490 ;
        RECT 76.945 156.210 77.225 156.490 ;
        RECT 77.345 156.210 77.625 156.490 ;
        RECT 77.745 156.210 78.025 156.490 ;
        RECT 79.845 153.490 80.125 153.770 ;
        RECT 80.245 153.490 80.525 153.770 ;
        RECT 80.645 153.490 80.925 153.770 ;
        RECT 81.045 153.490 81.325 153.770 ;
        RECT 76.545 150.770 76.825 151.050 ;
        RECT 76.945 150.770 77.225 151.050 ;
        RECT 77.345 150.770 77.625 151.050 ;
        RECT 77.745 150.770 78.025 151.050 ;
        RECT 88.620 188.850 88.900 189.130 ;
        RECT 89.020 188.850 89.300 189.130 ;
        RECT 89.420 188.850 89.700 189.130 ;
        RECT 89.820 188.850 90.100 189.130 ;
        RECT 91.920 186.130 92.200 186.410 ;
        RECT 92.320 186.130 92.600 186.410 ;
        RECT 92.720 186.130 93.000 186.410 ;
        RECT 93.120 186.130 93.400 186.410 ;
        RECT 100.695 188.850 100.975 189.130 ;
        RECT 101.095 188.850 101.375 189.130 ;
        RECT 101.495 188.850 101.775 189.130 ;
        RECT 101.895 188.850 102.175 189.130 ;
        RECT 88.620 183.410 88.900 183.690 ;
        RECT 89.020 183.410 89.300 183.690 ;
        RECT 89.420 183.410 89.700 183.690 ;
        RECT 89.820 183.410 90.100 183.690 ;
        RECT 91.920 180.690 92.200 180.970 ;
        RECT 92.320 180.690 92.600 180.970 ;
        RECT 92.720 180.690 93.000 180.970 ;
        RECT 93.120 180.690 93.400 180.970 ;
        RECT 88.620 177.970 88.900 178.250 ;
        RECT 89.020 177.970 89.300 178.250 ;
        RECT 89.420 177.970 89.700 178.250 ;
        RECT 89.820 177.970 90.100 178.250 ;
        RECT 91.920 175.250 92.200 175.530 ;
        RECT 92.320 175.250 92.600 175.530 ;
        RECT 92.720 175.250 93.000 175.530 ;
        RECT 93.120 175.250 93.400 175.530 ;
        RECT 103.995 191.570 104.275 191.850 ;
        RECT 104.395 191.570 104.675 191.850 ;
        RECT 104.795 191.570 105.075 191.850 ;
        RECT 105.195 191.570 105.475 191.850 ;
        RECT 103.995 186.130 104.275 186.410 ;
        RECT 104.395 186.130 104.675 186.410 ;
        RECT 104.795 186.130 105.075 186.410 ;
        RECT 105.195 186.130 105.475 186.410 ;
        RECT 116.070 191.570 116.350 191.850 ;
        RECT 116.470 191.570 116.750 191.850 ;
        RECT 116.870 191.570 117.150 191.850 ;
        RECT 117.270 191.570 117.550 191.850 ;
        RECT 100.695 183.410 100.975 183.690 ;
        RECT 101.095 183.410 101.375 183.690 ;
        RECT 101.495 183.410 101.775 183.690 ;
        RECT 101.895 183.410 102.175 183.690 ;
        RECT 88.620 172.530 88.900 172.810 ;
        RECT 89.020 172.530 89.300 172.810 ;
        RECT 89.420 172.530 89.700 172.810 ;
        RECT 89.820 172.530 90.100 172.810 ;
        RECT 20.405 149.825 20.705 150.125 ;
        RECT 49.415 147.950 49.895 148.430 ;
        RECT 79.845 148.050 80.125 148.330 ;
        RECT 80.245 148.050 80.525 148.330 ;
        RECT 80.645 148.050 80.925 148.330 ;
        RECT 81.045 148.050 81.325 148.330 ;
        RECT 19.630 147.565 19.960 147.865 ;
        RECT 25.545 143.440 26.260 144.195 ;
        RECT 21.070 142.980 21.370 143.280 ;
        RECT 86.060 154.510 86.340 154.790 ;
        RECT 91.920 169.810 92.200 170.090 ;
        RECT 92.320 169.810 92.600 170.090 ;
        RECT 92.720 169.810 93.000 170.090 ;
        RECT 93.120 169.810 93.400 170.090 ;
        RECT 100.695 177.970 100.975 178.250 ;
        RECT 101.095 177.970 101.375 178.250 ;
        RECT 101.495 177.970 101.775 178.250 ;
        RECT 101.895 177.970 102.175 178.250 ;
        RECT 100.695 172.530 100.975 172.810 ;
        RECT 101.095 172.530 101.375 172.810 ;
        RECT 101.495 172.530 101.775 172.810 ;
        RECT 101.895 172.530 102.175 172.810 ;
        RECT 88.620 167.090 88.900 167.370 ;
        RECT 89.020 167.090 89.300 167.370 ;
        RECT 89.420 167.090 89.700 167.370 ;
        RECT 89.820 167.090 90.100 167.370 ;
        RECT 88.620 161.650 88.900 161.930 ;
        RECT 89.020 161.650 89.300 161.930 ;
        RECT 89.420 161.650 89.700 161.930 ;
        RECT 89.820 161.650 90.100 161.930 ;
        RECT 91.920 164.370 92.200 164.650 ;
        RECT 92.320 164.370 92.600 164.650 ;
        RECT 92.720 164.370 93.000 164.650 ;
        RECT 93.120 164.370 93.400 164.650 ;
        RECT 91.920 158.930 92.200 159.210 ;
        RECT 92.320 158.930 92.600 159.210 ;
        RECT 92.720 158.930 93.000 159.210 ;
        RECT 93.120 158.930 93.400 159.210 ;
        RECT 88.620 156.210 88.900 156.490 ;
        RECT 89.020 156.210 89.300 156.490 ;
        RECT 89.420 156.210 89.700 156.490 ;
        RECT 89.820 156.210 90.100 156.490 ;
        RECT 91.920 153.490 92.200 153.770 ;
        RECT 92.320 153.490 92.600 153.770 ;
        RECT 92.720 153.490 93.000 153.770 ;
        RECT 93.120 153.490 93.400 153.770 ;
        RECT 100.695 167.090 100.975 167.370 ;
        RECT 101.095 167.090 101.375 167.370 ;
        RECT 101.495 167.090 101.775 167.370 ;
        RECT 101.895 167.090 102.175 167.370 ;
        RECT 100.695 161.650 100.975 161.930 ;
        RECT 101.095 161.650 101.375 161.930 ;
        RECT 101.495 161.650 101.775 161.930 ;
        RECT 101.895 161.650 102.175 161.930 ;
        RECT 103.995 180.690 104.275 180.970 ;
        RECT 104.395 180.690 104.675 180.970 ;
        RECT 104.795 180.690 105.075 180.970 ;
        RECT 105.195 180.690 105.475 180.970 ;
        RECT 103.995 175.250 104.275 175.530 ;
        RECT 104.395 175.250 104.675 175.530 ;
        RECT 104.795 175.250 105.075 175.530 ;
        RECT 105.195 175.250 105.475 175.530 ;
        RECT 103.995 169.810 104.275 170.090 ;
        RECT 104.395 169.810 104.675 170.090 ;
        RECT 104.795 169.810 105.075 170.090 ;
        RECT 105.195 169.810 105.475 170.090 ;
        RECT 103.995 164.370 104.275 164.650 ;
        RECT 104.395 164.370 104.675 164.650 ;
        RECT 104.795 164.370 105.075 164.650 ;
        RECT 105.195 164.370 105.475 164.650 ;
        RECT 100.695 156.210 100.975 156.490 ;
        RECT 101.095 156.210 101.375 156.490 ;
        RECT 101.495 156.210 101.775 156.490 ;
        RECT 101.895 156.210 102.175 156.490 ;
        RECT 88.620 150.770 88.900 151.050 ;
        RECT 89.020 150.770 89.300 151.050 ;
        RECT 89.420 150.770 89.700 151.050 ;
        RECT 89.820 150.770 90.100 151.050 ;
        RECT 103.995 158.930 104.275 159.210 ;
        RECT 104.395 158.930 104.675 159.210 ;
        RECT 104.795 158.930 105.075 159.210 ;
        RECT 105.195 158.930 105.475 159.210 ;
        RECT 103.995 153.490 104.275 153.770 ;
        RECT 104.395 153.490 104.675 153.770 ;
        RECT 104.795 153.490 105.075 153.770 ;
        RECT 105.195 153.490 105.475 153.770 ;
        RECT 100.695 150.770 100.975 151.050 ;
        RECT 101.095 150.770 101.375 151.050 ;
        RECT 101.495 150.770 101.775 151.050 ;
        RECT 101.895 150.770 102.175 151.050 ;
        RECT 120.100 189.190 120.380 189.470 ;
        RECT 112.770 188.850 113.050 189.130 ;
        RECT 113.170 188.850 113.450 189.130 ;
        RECT 113.570 188.850 113.850 189.130 ;
        RECT 113.970 188.850 114.250 189.130 ;
        RECT 116.070 186.130 116.350 186.410 ;
        RECT 116.470 186.130 116.750 186.410 ;
        RECT 116.870 186.130 117.150 186.410 ;
        RECT 117.270 186.130 117.550 186.410 ;
        RECT 112.770 183.410 113.050 183.690 ;
        RECT 113.170 183.410 113.450 183.690 ;
        RECT 113.570 183.410 113.850 183.690 ;
        RECT 113.970 183.410 114.250 183.690 ;
        RECT 112.770 177.970 113.050 178.250 ;
        RECT 113.170 177.970 113.450 178.250 ;
        RECT 113.570 177.970 113.850 178.250 ;
        RECT 113.970 177.970 114.250 178.250 ;
        RECT 116.070 180.690 116.350 180.970 ;
        RECT 116.470 180.690 116.750 180.970 ;
        RECT 116.870 180.690 117.150 180.970 ;
        RECT 117.270 180.690 117.550 180.970 ;
        RECT 112.770 172.530 113.050 172.810 ;
        RECT 113.170 172.530 113.450 172.810 ;
        RECT 113.570 172.530 113.850 172.810 ;
        RECT 113.970 172.530 114.250 172.810 ;
        RECT 112.770 167.090 113.050 167.370 ;
        RECT 113.170 167.090 113.450 167.370 ;
        RECT 113.570 167.090 113.850 167.370 ;
        RECT 113.970 167.090 114.250 167.370 ;
        RECT 116.070 175.250 116.350 175.530 ;
        RECT 116.470 175.250 116.750 175.530 ;
        RECT 116.870 175.250 117.150 175.530 ;
        RECT 117.270 175.250 117.550 175.530 ;
        RECT 116.070 169.810 116.350 170.090 ;
        RECT 116.470 169.810 116.750 170.090 ;
        RECT 116.870 169.810 117.150 170.090 ;
        RECT 117.270 169.810 117.550 170.090 ;
        RECT 112.770 161.650 113.050 161.930 ;
        RECT 113.170 161.650 113.450 161.930 ;
        RECT 113.570 161.650 113.850 161.930 ;
        RECT 113.970 161.650 114.250 161.930 ;
        RECT 116.070 164.370 116.350 164.650 ;
        RECT 116.470 164.370 116.750 164.650 ;
        RECT 116.870 164.370 117.150 164.650 ;
        RECT 117.270 164.370 117.550 164.650 ;
        RECT 116.070 158.930 116.350 159.210 ;
        RECT 116.470 158.930 116.750 159.210 ;
        RECT 116.870 158.930 117.150 159.210 ;
        RECT 117.270 158.930 117.550 159.210 ;
        RECT 112.770 156.210 113.050 156.490 ;
        RECT 113.170 156.210 113.450 156.490 ;
        RECT 113.570 156.210 113.850 156.490 ;
        RECT 113.970 156.210 114.250 156.490 ;
        RECT 116.070 153.490 116.350 153.770 ;
        RECT 116.470 153.490 116.750 153.770 ;
        RECT 116.870 153.490 117.150 153.770 ;
        RECT 117.270 153.490 117.550 153.770 ;
        RECT 112.770 150.770 113.050 151.050 ;
        RECT 113.170 150.770 113.450 151.050 ;
        RECT 113.570 150.770 113.850 151.050 ;
        RECT 113.970 150.770 114.250 151.050 ;
        RECT 120.100 153.830 120.380 154.110 ;
        RECT 91.920 148.050 92.200 148.330 ;
        RECT 92.320 148.050 92.600 148.330 ;
        RECT 92.720 148.050 93.000 148.330 ;
        RECT 93.120 148.050 93.400 148.330 ;
        RECT 103.995 148.050 104.275 148.330 ;
        RECT 104.395 148.050 104.675 148.330 ;
        RECT 104.795 148.050 105.075 148.330 ;
        RECT 105.195 148.050 105.475 148.330 ;
        RECT 116.070 148.050 116.350 148.330 ;
        RECT 116.470 148.050 116.750 148.330 ;
        RECT 116.870 148.050 117.150 148.330 ;
        RECT 117.270 148.050 117.550 148.330 ;
        RECT 80.300 139.095 81.150 139.945 ;
        RECT 110.375 139.260 110.885 139.820 ;
        RECT 88.155 135.325 88.705 135.875 ;
        RECT 152.060 135.300 152.660 135.900 ;
        RECT 13.070 123.935 13.935 124.915 ;
        RECT 46.565 121.910 46.865 122.210 ;
        RECT 20.185 111.855 20.485 112.155 ;
        RECT 19.410 109.595 19.740 109.895 ;
        RECT 1.365 82.730 2.055 83.240 ;
        RECT 103.640 109.010 103.930 109.290 ;
        RECT 25.325 105.470 26.040 106.225 ;
        RECT 20.850 105.010 21.150 105.310 ;
        RECT 44.585 88.970 44.885 89.270 ;
        RECT 49.350 88.610 50.010 89.310 ;
        RECT 88.130 101.815 88.730 102.415 ;
        RECT 103.540 101.980 103.890 102.290 ;
        RECT 42.855 75.775 43.250 76.125 ;
        RECT 42.860 73.480 43.255 73.830 ;
        RECT 1.320 62.900 1.940 63.690 ;
        RECT 32.960 71.970 33.340 72.280 ;
        RECT 27.570 69.705 27.905 70.030 ;
        RECT 49.470 68.890 50.090 69.680 ;
        RECT 27.470 67.450 27.770 67.740 ;
        RECT 34.540 64.690 34.850 64.970 ;
        RECT 27.730 63.340 28.065 63.665 ;
        RECT 53.395 61.225 53.760 61.605 ;
        RECT 28.780 59.195 29.190 59.545 ;
        RECT 34.220 59.225 34.670 59.575 ;
        RECT 23.180 56.600 23.630 57.180 ;
        RECT 23.630 48.930 25.220 50.170 ;
        RECT 1.280 35.295 2.220 36.155 ;
        RECT 55.655 56.860 56.090 57.345 ;
        RECT 101.265 88.800 101.545 89.080 ;
        RECT 101.665 88.800 101.945 89.080 ;
        RECT 102.065 88.800 102.345 89.080 ;
        RECT 102.465 88.800 102.745 89.080 ;
        RECT 116.560 88.800 116.840 89.080 ;
        RECT 116.960 88.800 117.240 89.080 ;
        RECT 117.360 88.800 117.640 89.080 ;
        RECT 117.760 88.800 118.040 89.080 ;
        RECT 131.855 88.800 132.135 89.080 ;
        RECT 132.255 88.800 132.535 89.080 ;
        RECT 132.655 88.800 132.935 89.080 ;
        RECT 133.055 88.800 133.335 89.080 ;
        RECT 151.870 89.140 152.150 89.420 ;
        RECT 147.150 88.800 147.430 89.080 ;
        RECT 147.550 88.800 147.830 89.080 ;
        RECT 147.950 88.800 148.230 89.080 ;
        RECT 148.350 88.800 148.630 89.080 ;
        RECT 97.965 86.080 98.245 86.360 ;
        RECT 98.365 86.080 98.645 86.360 ;
        RECT 98.765 86.080 99.045 86.360 ;
        RECT 99.165 86.080 99.445 86.360 ;
        RECT 101.265 83.360 101.545 83.640 ;
        RECT 101.665 83.360 101.945 83.640 ;
        RECT 102.065 83.360 102.345 83.640 ;
        RECT 102.465 83.360 102.745 83.640 ;
        RECT 97.965 80.640 98.245 80.920 ;
        RECT 98.365 80.640 98.645 80.920 ;
        RECT 98.765 80.640 99.045 80.920 ;
        RECT 99.165 80.640 99.445 80.920 ;
        RECT 105.870 79.620 106.150 79.900 ;
        RECT 101.265 77.920 101.545 78.200 ;
        RECT 101.665 77.920 101.945 78.200 ;
        RECT 102.065 77.920 102.345 78.200 ;
        RECT 102.465 77.920 102.745 78.200 ;
        RECT 97.965 75.200 98.245 75.480 ;
        RECT 98.365 75.200 98.645 75.480 ;
        RECT 98.765 75.200 99.045 75.480 ;
        RECT 99.165 75.200 99.445 75.480 ;
        RECT 101.265 72.480 101.545 72.760 ;
        RECT 101.665 72.480 101.945 72.760 ;
        RECT 102.065 72.480 102.345 72.760 ;
        RECT 102.465 72.480 102.745 72.760 ;
        RECT 97.965 69.760 98.245 70.040 ;
        RECT 98.365 69.760 98.645 70.040 ;
        RECT 98.765 69.760 99.045 70.040 ;
        RECT 99.165 69.760 99.445 70.040 ;
        RECT 101.265 67.040 101.545 67.320 ;
        RECT 101.665 67.040 101.945 67.320 ;
        RECT 102.065 67.040 102.345 67.320 ;
        RECT 102.465 67.040 102.745 67.320 ;
        RECT 97.965 64.320 98.245 64.600 ;
        RECT 98.365 64.320 98.645 64.600 ;
        RECT 98.765 64.320 99.045 64.600 ;
        RECT 99.165 64.320 99.445 64.600 ;
        RECT 101.265 61.600 101.545 61.880 ;
        RECT 101.665 61.600 101.945 61.880 ;
        RECT 102.065 61.600 102.345 61.880 ;
        RECT 102.465 61.600 102.745 61.880 ;
        RECT 88.155 38.685 88.705 39.235 ;
        RECT 90.230 38.820 90.510 39.100 ;
        RECT 97.965 58.880 98.245 59.160 ;
        RECT 98.365 58.880 98.645 59.160 ;
        RECT 98.765 58.880 99.045 59.160 ;
        RECT 99.165 58.880 99.445 59.160 ;
        RECT 101.265 56.160 101.545 56.440 ;
        RECT 101.665 56.160 101.945 56.440 ;
        RECT 102.065 56.160 102.345 56.440 ;
        RECT 102.465 56.160 102.745 56.440 ;
        RECT 97.965 53.440 98.245 53.720 ;
        RECT 98.365 53.440 98.645 53.720 ;
        RECT 98.765 53.440 99.045 53.720 ;
        RECT 99.165 53.440 99.445 53.720 ;
        RECT 97.965 48.000 98.245 48.280 ;
        RECT 98.365 48.000 98.645 48.280 ;
        RECT 98.765 48.000 99.045 48.280 ;
        RECT 99.165 48.000 99.445 48.280 ;
        RECT 97.965 42.560 98.245 42.840 ;
        RECT 98.365 42.560 98.645 42.840 ;
        RECT 98.765 42.560 99.045 42.840 ;
        RECT 99.165 42.560 99.445 42.840 ;
        RECT 98.970 38.140 99.250 38.420 ;
        RECT 101.265 50.720 101.545 51.000 ;
        RECT 101.665 50.720 101.945 51.000 ;
        RECT 102.065 50.720 102.345 51.000 ;
        RECT 102.465 50.720 102.745 51.000 ;
        RECT 101.265 45.280 101.545 45.560 ;
        RECT 101.665 45.280 101.945 45.560 ;
        RECT 102.065 45.280 102.345 45.560 ;
        RECT 102.465 45.280 102.745 45.560 ;
        RECT 101.265 39.840 101.545 40.120 ;
        RECT 101.665 39.840 101.945 40.120 ;
        RECT 102.065 39.840 102.345 40.120 ;
        RECT 102.465 39.840 102.745 40.120 ;
        RECT 97.965 37.120 98.245 37.400 ;
        RECT 98.365 37.120 98.645 37.400 ;
        RECT 98.765 37.120 99.045 37.400 ;
        RECT 99.165 37.120 99.445 37.400 ;
        RECT 101.265 34.400 101.545 34.680 ;
        RECT 101.665 34.400 101.945 34.680 ;
        RECT 102.065 34.400 102.345 34.680 ;
        RECT 102.465 34.400 102.745 34.680 ;
        RECT 97.965 31.680 98.245 31.960 ;
        RECT 98.365 31.680 98.645 31.960 ;
        RECT 98.765 31.680 99.045 31.960 ;
        RECT 99.165 31.680 99.445 31.960 ;
        RECT 113.260 86.080 113.540 86.360 ;
        RECT 113.660 86.080 113.940 86.360 ;
        RECT 114.060 86.080 114.340 86.360 ;
        RECT 114.460 86.080 114.740 86.360 ;
        RECT 128.555 86.080 128.835 86.360 ;
        RECT 128.955 86.080 129.235 86.360 ;
        RECT 129.355 86.080 129.635 86.360 ;
        RECT 129.755 86.080 130.035 86.360 ;
        RECT 116.560 83.360 116.840 83.640 ;
        RECT 116.960 83.360 117.240 83.640 ;
        RECT 117.360 83.360 117.640 83.640 ;
        RECT 117.760 83.360 118.040 83.640 ;
        RECT 113.260 80.640 113.540 80.920 ;
        RECT 113.660 80.640 113.940 80.920 ;
        RECT 114.060 80.640 114.340 80.920 ;
        RECT 114.460 80.640 114.740 80.920 ;
        RECT 116.560 77.920 116.840 78.200 ;
        RECT 116.960 77.920 117.240 78.200 ;
        RECT 117.360 77.920 117.640 78.200 ;
        RECT 117.760 77.920 118.040 78.200 ;
        RECT 113.260 75.200 113.540 75.480 ;
        RECT 113.660 75.200 113.940 75.480 ;
        RECT 114.060 75.200 114.340 75.480 ;
        RECT 114.460 75.200 114.740 75.480 ;
        RECT 113.260 69.760 113.540 70.040 ;
        RECT 113.660 69.760 113.940 70.040 ;
        RECT 114.060 69.760 114.340 70.040 ;
        RECT 114.460 69.760 114.740 70.040 ;
        RECT 113.260 64.320 113.540 64.600 ;
        RECT 113.660 64.320 113.940 64.600 ;
        RECT 114.060 64.320 114.340 64.600 ;
        RECT 114.460 64.320 114.740 64.600 ;
        RECT 116.560 72.480 116.840 72.760 ;
        RECT 116.960 72.480 117.240 72.760 ;
        RECT 117.360 72.480 117.640 72.760 ;
        RECT 117.760 72.480 118.040 72.760 ;
        RECT 116.560 67.040 116.840 67.320 ;
        RECT 116.960 67.040 117.240 67.320 ;
        RECT 117.360 67.040 117.640 67.320 ;
        RECT 117.760 67.040 118.040 67.320 ;
        RECT 131.855 83.360 132.135 83.640 ;
        RECT 132.255 83.360 132.535 83.640 ;
        RECT 132.655 83.360 132.935 83.640 ;
        RECT 133.055 83.360 133.335 83.640 ;
        RECT 128.555 80.640 128.835 80.920 ;
        RECT 128.955 80.640 129.235 80.920 ;
        RECT 129.355 80.640 129.635 80.920 ;
        RECT 129.755 80.640 130.035 80.920 ;
        RECT 127.490 78.940 127.770 79.220 ;
        RECT 128.555 75.200 128.835 75.480 ;
        RECT 128.955 75.200 129.235 75.480 ;
        RECT 129.355 75.200 129.635 75.480 ;
        RECT 129.755 75.200 130.035 75.480 ;
        RECT 133.930 78.260 134.210 78.540 ;
        RECT 131.855 77.920 132.135 78.200 ;
        RECT 132.255 77.920 132.535 78.200 ;
        RECT 132.655 77.920 132.935 78.200 ;
        RECT 133.055 77.920 133.335 78.200 ;
        RECT 136.230 78.260 136.510 78.540 ;
        RECT 143.850 86.080 144.130 86.360 ;
        RECT 144.250 86.080 144.530 86.360 ;
        RECT 144.650 86.080 144.930 86.360 ;
        RECT 145.050 86.080 145.330 86.360 ;
        RECT 143.850 80.640 144.130 80.920 ;
        RECT 144.250 80.640 144.530 80.920 ;
        RECT 144.650 80.640 144.930 80.920 ;
        RECT 145.050 80.640 145.330 80.920 ;
        RECT 147.150 83.360 147.430 83.640 ;
        RECT 147.550 83.360 147.830 83.640 ;
        RECT 147.950 83.360 148.230 83.640 ;
        RECT 148.350 83.360 148.630 83.640 ;
        RECT 131.855 72.480 132.135 72.760 ;
        RECT 132.255 72.480 132.535 72.760 ;
        RECT 132.655 72.480 132.935 72.760 ;
        RECT 133.055 72.480 133.335 72.760 ;
        RECT 116.560 61.600 116.840 61.880 ;
        RECT 116.960 61.600 117.240 61.880 ;
        RECT 117.360 61.600 117.640 61.880 ;
        RECT 117.760 61.600 118.040 61.880 ;
        RECT 113.260 58.880 113.540 59.160 ;
        RECT 113.660 58.880 113.940 59.160 ;
        RECT 114.060 58.880 114.340 59.160 ;
        RECT 114.460 58.880 114.740 59.160 ;
        RECT 116.560 56.160 116.840 56.440 ;
        RECT 116.960 56.160 117.240 56.440 ;
        RECT 117.360 56.160 117.640 56.440 ;
        RECT 117.760 56.160 118.040 56.440 ;
        RECT 113.260 53.440 113.540 53.720 ;
        RECT 113.660 53.440 113.940 53.720 ;
        RECT 114.060 53.440 114.340 53.720 ;
        RECT 114.460 53.440 114.740 53.720 ;
        RECT 116.560 50.720 116.840 51.000 ;
        RECT 116.960 50.720 117.240 51.000 ;
        RECT 117.360 50.720 117.640 51.000 ;
        RECT 117.760 50.720 118.040 51.000 ;
        RECT 113.260 48.000 113.540 48.280 ;
        RECT 113.660 48.000 113.940 48.280 ;
        RECT 114.060 48.000 114.340 48.280 ;
        RECT 114.460 48.000 114.740 48.280 ;
        RECT 116.560 45.280 116.840 45.560 ;
        RECT 116.960 45.280 117.240 45.560 ;
        RECT 117.360 45.280 117.640 45.560 ;
        RECT 117.760 45.280 118.040 45.560 ;
        RECT 113.260 42.560 113.540 42.840 ;
        RECT 113.660 42.560 113.940 42.840 ;
        RECT 114.060 42.560 114.340 42.840 ;
        RECT 114.460 42.560 114.740 42.840 ;
        RECT 116.560 39.840 116.840 40.120 ;
        RECT 116.960 39.840 117.240 40.120 ;
        RECT 117.360 39.840 117.640 40.120 ;
        RECT 117.760 39.840 118.040 40.120 ;
        RECT 128.555 69.760 128.835 70.040 ;
        RECT 128.955 69.760 129.235 70.040 ;
        RECT 129.355 69.760 129.635 70.040 ;
        RECT 129.755 69.760 130.035 70.040 ;
        RECT 131.855 67.040 132.135 67.320 ;
        RECT 132.255 67.040 132.535 67.320 ;
        RECT 132.655 67.040 132.935 67.320 ;
        RECT 133.055 67.040 133.335 67.320 ;
        RECT 140.830 78.940 141.110 79.220 ;
        RECT 143.850 75.200 144.130 75.480 ;
        RECT 144.250 75.200 144.530 75.480 ;
        RECT 144.650 75.200 144.930 75.480 ;
        RECT 145.050 75.200 145.330 75.480 ;
        RECT 147.150 77.920 147.430 78.200 ;
        RECT 147.550 77.920 147.830 78.200 ;
        RECT 147.950 77.920 148.230 78.200 ;
        RECT 148.350 77.920 148.630 78.200 ;
        RECT 143.850 69.760 144.130 70.040 ;
        RECT 144.250 69.760 144.530 70.040 ;
        RECT 144.650 69.760 144.930 70.040 ;
        RECT 145.050 69.760 145.330 70.040 ;
        RECT 147.150 72.480 147.430 72.760 ;
        RECT 147.550 72.480 147.830 72.760 ;
        RECT 147.950 72.480 148.230 72.760 ;
        RECT 148.350 72.480 148.630 72.760 ;
        RECT 128.555 64.320 128.835 64.600 ;
        RECT 128.955 64.320 129.235 64.600 ;
        RECT 129.355 64.320 129.635 64.600 ;
        RECT 129.755 64.320 130.035 64.600 ;
        RECT 131.855 61.600 132.135 61.880 ;
        RECT 132.255 61.600 132.535 61.880 ;
        RECT 132.655 61.600 132.935 61.880 ;
        RECT 133.055 61.600 133.335 61.880 ;
        RECT 143.850 64.320 144.130 64.600 ;
        RECT 144.250 64.320 144.530 64.600 ;
        RECT 144.650 64.320 144.930 64.600 ;
        RECT 145.050 64.320 145.330 64.600 ;
        RECT 128.555 58.880 128.835 59.160 ;
        RECT 128.955 58.880 129.235 59.160 ;
        RECT 129.355 58.880 129.635 59.160 ;
        RECT 129.755 58.880 130.035 59.160 ;
        RECT 143.850 58.880 144.130 59.160 ;
        RECT 144.250 58.880 144.530 59.160 ;
        RECT 144.650 58.880 144.930 59.160 ;
        RECT 145.050 58.880 145.330 59.160 ;
        RECT 128.555 53.440 128.835 53.720 ;
        RECT 128.955 53.440 129.235 53.720 ;
        RECT 129.355 53.440 129.635 53.720 ;
        RECT 129.755 53.440 130.035 53.720 ;
        RECT 131.855 56.160 132.135 56.440 ;
        RECT 132.255 56.160 132.535 56.440 ;
        RECT 132.655 56.160 132.935 56.440 ;
        RECT 133.055 56.160 133.335 56.440 ;
        RECT 128.555 48.000 128.835 48.280 ;
        RECT 128.955 48.000 129.235 48.280 ;
        RECT 129.355 48.000 129.635 48.280 ;
        RECT 129.755 48.000 130.035 48.280 ;
        RECT 131.855 50.720 132.135 51.000 ;
        RECT 132.255 50.720 132.535 51.000 ;
        RECT 132.655 50.720 132.935 51.000 ;
        RECT 133.055 50.720 133.335 51.000 ;
        RECT 131.855 45.280 132.135 45.560 ;
        RECT 132.255 45.280 132.535 45.560 ;
        RECT 132.655 45.280 132.935 45.560 ;
        RECT 133.055 45.280 133.335 45.560 ;
        RECT 112.770 38.140 113.050 38.420 ;
        RECT 113.260 37.120 113.540 37.400 ;
        RECT 113.660 37.120 113.940 37.400 ;
        RECT 114.060 37.120 114.340 37.400 ;
        RECT 114.460 37.120 114.740 37.400 ;
        RECT 117.830 37.460 118.110 37.740 ;
        RECT 116.560 34.400 116.840 34.680 ;
        RECT 116.960 34.400 117.240 34.680 ;
        RECT 117.360 34.400 117.640 34.680 ;
        RECT 117.760 34.400 118.040 34.680 ;
        RECT 121.510 35.420 121.790 35.700 ;
        RECT 113.260 31.680 113.540 31.960 ;
        RECT 113.660 31.680 113.940 31.960 ;
        RECT 114.060 31.680 114.340 31.960 ;
        RECT 114.460 31.680 114.740 31.960 ;
        RECT 128.555 42.560 128.835 42.840 ;
        RECT 128.955 42.560 129.235 42.840 ;
        RECT 129.355 42.560 129.635 42.840 ;
        RECT 129.755 42.560 130.035 42.840 ;
        RECT 131.855 39.840 132.135 40.120 ;
        RECT 132.255 39.840 132.535 40.120 ;
        RECT 132.655 39.840 132.935 40.120 ;
        RECT 133.055 39.840 133.335 40.120 ;
        RECT 143.850 53.440 144.130 53.720 ;
        RECT 144.250 53.440 144.530 53.720 ;
        RECT 144.650 53.440 144.930 53.720 ;
        RECT 145.050 53.440 145.330 53.720 ;
        RECT 150.490 68.740 150.770 69.020 ;
        RECT 147.150 67.040 147.430 67.320 ;
        RECT 147.550 67.040 147.830 67.320 ;
        RECT 147.950 67.040 148.230 67.320 ;
        RECT 148.350 67.040 148.630 67.320 ;
        RECT 147.150 61.600 147.430 61.880 ;
        RECT 147.550 61.600 147.830 61.880 ;
        RECT 147.950 61.600 148.230 61.880 ;
        RECT 148.350 61.600 148.630 61.880 ;
        RECT 147.150 56.160 147.430 56.440 ;
        RECT 147.550 56.160 147.830 56.440 ;
        RECT 147.950 56.160 148.230 56.440 ;
        RECT 148.350 56.160 148.630 56.440 ;
        RECT 147.150 50.720 147.430 51.000 ;
        RECT 147.550 50.720 147.830 51.000 ;
        RECT 147.950 50.720 148.230 51.000 ;
        RECT 148.350 50.720 148.630 51.000 ;
        RECT 150.490 48.340 150.770 48.620 ;
        RECT 143.850 48.000 144.130 48.280 ;
        RECT 144.250 48.000 144.530 48.280 ;
        RECT 144.650 48.000 144.930 48.280 ;
        RECT 145.050 48.000 145.330 48.280 ;
        RECT 147.150 45.280 147.430 45.560 ;
        RECT 147.550 45.280 147.830 45.560 ;
        RECT 147.950 45.280 148.230 45.560 ;
        RECT 148.350 45.280 148.630 45.560 ;
        RECT 127.030 37.460 127.310 37.740 ;
        RECT 128.555 37.120 128.835 37.400 ;
        RECT 128.955 37.120 129.235 37.400 ;
        RECT 129.355 37.120 129.635 37.400 ;
        RECT 129.755 37.120 130.035 37.400 ;
        RECT 127.030 35.420 127.310 35.700 ;
        RECT 131.855 34.400 132.135 34.680 ;
        RECT 132.255 34.400 132.535 34.680 ;
        RECT 132.655 34.400 132.935 34.680 ;
        RECT 133.055 34.400 133.335 34.680 ;
        RECT 143.850 42.560 144.130 42.840 ;
        RECT 144.250 42.560 144.530 42.840 ;
        RECT 144.650 42.560 144.930 42.840 ;
        RECT 145.050 42.560 145.330 42.840 ;
        RECT 147.150 39.840 147.430 40.120 ;
        RECT 147.550 39.840 147.830 40.120 ;
        RECT 147.950 39.840 148.230 40.120 ;
        RECT 148.350 39.840 148.630 40.120 ;
        RECT 143.850 37.120 144.130 37.400 ;
        RECT 144.250 37.120 144.530 37.400 ;
        RECT 144.650 37.120 144.930 37.400 ;
        RECT 145.050 37.120 145.330 37.400 ;
        RECT 128.555 31.680 128.835 31.960 ;
        RECT 128.955 31.680 129.235 31.960 ;
        RECT 129.355 31.680 129.635 31.960 ;
        RECT 129.755 31.680 130.035 31.960 ;
        RECT 147.150 34.400 147.430 34.680 ;
        RECT 147.550 34.400 147.830 34.680 ;
        RECT 147.950 34.400 148.230 34.680 ;
        RECT 148.350 34.400 148.630 34.680 ;
        RECT 143.850 31.680 144.130 31.960 ;
        RECT 144.250 31.680 144.530 31.960 ;
        RECT 144.650 31.680 144.930 31.960 ;
        RECT 145.050 31.680 145.330 31.960 ;
        RECT 1.280 23.810 2.220 24.670 ;
        RECT 101.265 28.960 101.545 29.240 ;
        RECT 101.665 28.960 101.945 29.240 ;
        RECT 102.065 28.960 102.345 29.240 ;
        RECT 102.465 28.960 102.745 29.240 ;
        RECT 116.560 28.960 116.840 29.240 ;
        RECT 116.960 28.960 117.240 29.240 ;
        RECT 117.360 28.960 117.640 29.240 ;
        RECT 117.760 28.960 118.040 29.240 ;
        RECT 131.855 28.960 132.135 29.240 ;
        RECT 132.255 28.960 132.535 29.240 ;
        RECT 132.655 28.960 132.935 29.240 ;
        RECT 133.055 28.960 133.335 29.240 ;
        RECT 147.150 28.960 147.430 29.240 ;
        RECT 147.550 28.960 147.830 29.240 ;
        RECT 147.950 28.960 148.230 29.240 ;
        RECT 148.350 28.960 148.630 29.240 ;
        RECT 151.870 27.940 152.150 28.220 ;
        RECT 59.095 20.600 59.375 20.880 ;
        RECT 8.560 16.620 9.610 17.985 ;
        RECT 71.345 15.365 71.645 15.665 ;
        RECT 69.885 14.660 70.185 14.960 ;
        RECT 68.680 13.750 68.980 14.050 ;
        RECT 67.725 13.090 68.025 13.390 ;
        RECT 66.770 12.500 67.070 12.800 ;
        RECT 65.745 11.700 66.045 12.000 ;
        RECT 64.760 10.955 65.060 11.255 ;
        RECT 63.760 9.880 64.060 10.180 ;
        RECT 62.540 9.110 62.840 9.410 ;
        RECT 53.335 8.005 53.805 8.460 ;
        RECT 24.180 6.915 24.550 7.270 ;
        RECT 83.210 7.760 83.645 8.180 ;
      LAYER met3 ;
        RECT 84.840 222.455 85.360 222.940 ;
        RECT 88.500 222.470 89.020 222.955 ;
        RECT 154.280 222.745 156.080 224.045 ;
        RECT 66.565 220.465 66.885 220.845 ;
        RECT 70.205 220.505 70.525 220.885 ;
        RECT 147.325 220.800 147.975 221.480 ;
        RECT 46.525 219.215 46.905 219.225 ;
        RECT 66.575 219.215 66.875 220.465 ;
        RECT 46.525 218.915 66.875 219.215 ;
        RECT 46.525 218.905 46.905 218.915 ;
        RECT 44.545 217.925 44.925 217.935 ;
        RECT 70.215 217.925 70.515 220.505 ;
        RECT 143.605 218.905 144.325 219.620 ;
        RECT 44.545 217.625 70.515 217.925 ;
        RECT 44.545 217.615 44.925 217.625 ;
        RECT 139.920 216.725 140.640 217.440 ;
        RECT 153.605 216.750 154.255 217.405 ;
        RECT 136.265 215.055 136.985 215.770 ;
        RECT 153.840 215.090 154.490 215.745 ;
        RECT 4.105 213.605 4.550 213.665 ;
        RECT 62.775 213.605 63.355 213.670 ;
        RECT 4.105 213.290 63.355 213.605 ;
        RECT 4.105 213.265 4.550 213.290 ;
        RECT 62.775 213.235 63.355 213.290 ;
        RECT 4.955 211.330 5.675 211.770 ;
        RECT 3.475 207.405 4.045 207.825 ;
        RECT 1.005 193.685 2.505 195.185 ;
        RECT 1.000 82.525 2.500 83.410 ;
        RECT 3.565 66.105 3.870 207.405 ;
        RECT 5.055 73.575 5.425 211.330 ;
        RECT 154.820 210.275 155.425 222.745 ;
        RECT 157.225 221.420 157.825 221.425 ;
        RECT 157.200 220.830 157.850 221.420 ;
        RECT 157.225 220.825 157.825 220.830 ;
        RECT 155.965 219.555 156.615 219.590 ;
        RECT 155.955 218.965 156.615 219.555 ;
        RECT 155.965 218.935 156.615 218.965 ;
        RECT 54.615 209.670 155.425 210.275 ;
        RECT 14.200 159.815 41.495 160.795 ;
        RECT 14.200 125.235 15.180 159.815 ;
        RECT 31.815 153.265 35.675 155.665 ;
        RECT 20.320 149.735 20.845 150.215 ;
        RECT 19.600 147.855 20.050 147.925 ;
        RECT 23.980 147.855 26.380 149.700 ;
        RECT 31.815 149.665 35.675 152.065 ;
        RECT 19.600 147.555 26.380 147.855 ;
        RECT 19.600 147.505 20.050 147.555 ;
        RECT 23.980 145.840 26.380 147.555 ;
        RECT 31.815 146.065 35.675 148.465 ;
        RECT 20.915 142.840 21.550 143.395 ;
        RECT 25.335 143.245 26.440 144.355 ;
        RECT 31.815 142.465 35.675 144.865 ;
        RECT 31.815 138.865 35.675 141.265 ;
        RECT 31.815 135.265 35.675 137.665 ;
        RECT 31.815 131.665 35.675 134.065 ;
        RECT 31.815 128.065 35.675 130.465 ;
        RECT 12.350 123.940 15.180 125.235 ;
        RECT 31.815 124.465 35.675 126.865 ;
        RECT 40.515 125.430 41.495 159.815 ;
        RECT 54.615 154.275 55.220 209.670 ;
        RECT 76.495 194.265 78.075 194.595 ;
        RECT 88.570 194.265 90.150 194.595 ;
        RECT 100.645 194.265 102.225 194.595 ;
        RECT 112.720 194.265 114.300 194.595 ;
        RECT 79.795 191.545 81.375 191.875 ;
        RECT 91.870 191.545 93.450 191.875 ;
        RECT 103.945 191.545 105.525 191.875 ;
        RECT 116.020 191.545 117.600 191.875 ;
        RECT 65.730 189.480 69.730 189.630 ;
        RECT 70.395 189.480 70.725 189.495 ;
        RECT 65.730 189.180 70.725 189.480 ;
        RECT 65.730 189.030 69.730 189.180 ;
        RECT 70.395 189.165 70.725 189.180 ;
        RECT 120.075 189.480 120.405 189.495 ;
        RECT 121.500 189.480 129.575 189.630 ;
        RECT 120.075 189.180 129.575 189.480 ;
        RECT 120.075 189.165 120.405 189.180 ;
        RECT 76.495 188.825 78.075 189.155 ;
        RECT 88.570 188.825 90.150 189.155 ;
        RECT 100.645 188.825 102.225 189.155 ;
        RECT 112.720 188.825 114.300 189.155 ;
        RECT 121.500 189.030 129.575 189.180 ;
        RECT 79.795 186.105 81.375 186.435 ;
        RECT 91.870 186.105 93.450 186.435 ;
        RECT 103.945 186.105 105.525 186.435 ;
        RECT 116.020 186.105 117.600 186.435 ;
        RECT 76.495 183.385 78.075 183.715 ;
        RECT 88.570 183.385 90.150 183.715 ;
        RECT 100.645 183.385 102.225 183.715 ;
        RECT 112.720 183.385 114.300 183.715 ;
        RECT 79.795 180.665 81.375 180.995 ;
        RECT 91.870 180.665 93.450 180.995 ;
        RECT 103.945 180.665 105.525 180.995 ;
        RECT 116.020 180.665 117.600 180.995 ;
        RECT 76.495 177.945 78.075 178.275 ;
        RECT 88.570 177.945 90.150 178.275 ;
        RECT 100.645 177.945 102.225 178.275 ;
        RECT 112.720 177.945 114.300 178.275 ;
        RECT 79.795 175.225 81.375 175.555 ;
        RECT 91.870 175.225 93.450 175.555 ;
        RECT 103.945 175.225 105.525 175.555 ;
        RECT 116.020 175.225 117.600 175.555 ;
        RECT 76.495 172.505 78.075 172.835 ;
        RECT 88.570 172.505 90.150 172.835 ;
        RECT 100.645 172.505 102.225 172.835 ;
        RECT 112.720 172.505 114.300 172.835 ;
        RECT 79.795 169.785 81.375 170.115 ;
        RECT 91.870 169.785 93.450 170.115 ;
        RECT 103.945 169.785 105.525 170.115 ;
        RECT 116.020 169.785 117.600 170.115 ;
        RECT 76.495 167.065 78.075 167.395 ;
        RECT 88.570 167.065 90.150 167.395 ;
        RECT 100.645 167.065 102.225 167.395 ;
        RECT 112.720 167.065 114.300 167.395 ;
        RECT 79.795 164.345 81.375 164.675 ;
        RECT 91.870 164.345 93.450 164.675 ;
        RECT 103.945 164.345 105.525 164.675 ;
        RECT 116.020 164.345 117.600 164.675 ;
        RECT 76.495 161.625 78.075 161.955 ;
        RECT 88.570 161.625 90.150 161.955 ;
        RECT 100.645 161.625 102.225 161.955 ;
        RECT 112.720 161.625 114.300 161.955 ;
        RECT 79.795 158.905 81.375 159.235 ;
        RECT 91.870 158.905 93.450 159.235 ;
        RECT 103.945 158.905 105.525 159.235 ;
        RECT 116.020 158.905 117.600 159.235 ;
        RECT 76.495 156.185 78.075 156.515 ;
        RECT 88.570 156.185 90.150 156.515 ;
        RECT 100.645 156.185 102.225 156.515 ;
        RECT 112.720 156.185 114.300 156.515 ;
        RECT 86.035 154.800 86.365 154.815 ;
        RECT 78.920 154.500 86.365 154.800 ;
        RECT 54.615 154.270 66.305 154.275 ;
        RECT 54.615 154.120 69.730 154.270 ;
        RECT 78.920 154.120 79.220 154.500 ;
        RECT 86.035 154.485 86.365 154.500 ;
        RECT 54.615 153.820 79.220 154.120 ;
        RECT 120.075 154.120 120.405 154.135 ;
        RECT 121.500 154.120 133.170 154.270 ;
        RECT 120.075 153.820 133.170 154.120 ;
        RECT 54.615 153.670 69.730 153.820 ;
        RECT 120.075 153.805 120.405 153.820 ;
        RECT 49.000 147.760 50.500 148.755 ;
        RECT 64.990 128.510 65.590 153.670 ;
        RECT 79.795 153.465 81.375 153.795 ;
        RECT 91.870 153.465 93.450 153.795 ;
        RECT 103.945 153.465 105.525 153.795 ;
        RECT 116.020 153.465 117.600 153.795 ;
        RECT 121.500 153.670 133.170 153.820 ;
        RECT 76.495 150.745 78.075 151.075 ;
        RECT 88.570 150.745 90.150 151.075 ;
        RECT 100.645 150.745 102.225 151.075 ;
        RECT 112.720 150.745 114.300 151.075 ;
        RECT 79.795 148.025 81.375 148.355 ;
        RECT 91.870 148.025 93.450 148.355 ;
        RECT 103.945 148.025 105.525 148.355 ;
        RECT 116.020 148.025 117.600 148.355 ;
        RECT 80.195 138.950 81.260 140.035 ;
        RECT 110.180 139.050 111.080 139.950 ;
        RECT 64.990 127.910 83.550 128.510 ;
        RECT 78.590 125.430 80.430 125.685 ;
        RECT 12.350 123.435 14.535 123.940 ;
        RECT 34.270 122.855 34.690 124.465 ;
        RECT 40.515 124.450 80.430 125.430 ;
        RECT 78.590 124.050 80.430 124.450 ;
        RECT 34.270 122.435 40.695 122.855 ;
        RECT 31.595 115.295 35.455 117.695 ;
        RECT 20.100 111.765 20.625 112.245 ;
        RECT 19.380 109.885 19.830 109.955 ;
        RECT 23.760 109.885 26.160 111.730 ;
        RECT 31.595 111.695 35.455 114.095 ;
        RECT 19.380 109.585 26.160 109.885 ;
        RECT 19.380 109.535 19.830 109.585 ;
        RECT 23.760 107.870 26.160 109.585 ;
        RECT 31.595 108.095 35.455 110.495 ;
        RECT 20.695 104.870 21.330 105.425 ;
        RECT 25.115 105.275 26.220 106.385 ;
        RECT 31.595 104.495 35.455 106.895 ;
        RECT 31.595 100.895 35.455 103.295 ;
        RECT 31.595 97.295 35.455 99.695 ;
        RECT 31.595 93.695 35.455 96.095 ;
        RECT 31.595 90.095 35.455 92.495 ;
        RECT 31.595 86.495 35.455 88.895 ;
        RECT 33.980 73.780 34.360 86.495 ;
        RECT 40.125 76.210 40.545 122.435 ;
        RECT 46.315 121.625 47.120 122.425 ;
        RECT 44.310 88.715 45.115 89.515 ;
        RECT 49.000 88.350 50.500 89.630 ;
        RECT 82.950 80.060 83.550 127.910 ;
        RECT 88.130 102.440 88.730 135.900 ;
        RECT 152.035 135.245 152.685 135.925 ;
        RECT 103.490 108.900 104.040 109.320 ;
        RECT 103.620 102.460 103.970 108.900 ;
        RECT 88.105 101.790 88.755 102.440 ;
        RECT 103.270 101.850 104.190 102.460 ;
        RECT 151.845 89.430 152.175 89.445 ;
        RECT 153.825 89.430 157.825 89.580 ;
        RECT 151.845 89.130 157.825 89.430 ;
        RECT 151.845 89.115 152.175 89.130 ;
        RECT 101.215 88.775 102.795 89.105 ;
        RECT 116.510 88.775 118.090 89.105 ;
        RECT 131.805 88.775 133.385 89.105 ;
        RECT 147.100 88.775 148.680 89.105 ;
        RECT 153.825 88.980 157.825 89.130 ;
        RECT 97.915 86.055 99.495 86.385 ;
        RECT 113.210 86.055 114.790 86.385 ;
        RECT 128.505 86.055 130.085 86.385 ;
        RECT 143.800 86.055 145.380 86.385 ;
        RECT 101.215 83.335 102.795 83.665 ;
        RECT 116.510 83.335 118.090 83.665 ;
        RECT 131.805 83.335 133.385 83.665 ;
        RECT 147.100 83.335 148.680 83.665 ;
        RECT 97.915 80.615 99.495 80.945 ;
        RECT 113.210 80.615 114.790 80.945 ;
        RECT 128.505 80.615 130.085 80.945 ;
        RECT 143.800 80.615 145.380 80.945 ;
        RECT 82.950 79.910 89.540 80.060 ;
        RECT 105.845 79.910 106.175 79.925 ;
        RECT 82.950 79.610 106.175 79.910 ;
        RECT 82.950 79.460 89.540 79.610 ;
        RECT 105.845 79.595 106.175 79.610 ;
        RECT 127.465 79.230 127.795 79.245 ;
        RECT 140.805 79.230 141.135 79.245 ;
        RECT 127.465 78.930 141.135 79.230 ;
        RECT 127.465 78.915 127.795 78.930 ;
        RECT 140.805 78.915 141.135 78.930 ;
        RECT 133.905 78.550 134.235 78.565 ;
        RECT 136.205 78.550 136.535 78.565 ;
        RECT 133.905 78.250 136.535 78.550 ;
        RECT 133.905 78.235 134.235 78.250 ;
        RECT 136.205 78.235 136.535 78.250 ;
        RECT 101.215 77.895 102.795 78.225 ;
        RECT 116.510 77.895 118.090 78.225 ;
        RECT 131.805 77.895 133.385 78.225 ;
        RECT 147.100 77.895 148.680 78.225 ;
        RECT 42.615 76.210 43.490 76.380 ;
        RECT 40.125 75.790 43.490 76.210 ;
        RECT 42.615 75.545 43.490 75.790 ;
        RECT 97.915 75.175 99.495 75.505 ;
        RECT 113.210 75.175 114.790 75.505 ;
        RECT 128.505 75.175 130.085 75.505 ;
        RECT 143.800 75.175 145.380 75.505 ;
        RECT 42.625 73.780 43.500 74.150 ;
        RECT 5.055 73.205 33.330 73.575 ;
        RECT 33.980 73.400 43.500 73.780 ;
        RECT 32.960 72.650 33.330 73.205 ;
        RECT 42.625 73.115 43.500 73.400 ;
        RECT 32.960 72.475 33.340 72.650 ;
        RECT 32.795 71.800 33.470 72.475 ;
        RECT 101.215 72.455 102.795 72.785 ;
        RECT 116.510 72.455 118.090 72.785 ;
        RECT 131.805 72.455 133.385 72.785 ;
        RECT 147.100 72.455 148.680 72.785 ;
        RECT 27.400 69.580 28.085 70.140 ;
        RECT 48.990 68.440 50.510 70.220 ;
        RECT 97.915 69.735 99.495 70.065 ;
        RECT 113.210 69.735 114.790 70.065 ;
        RECT 128.505 69.735 130.085 70.065 ;
        RECT 143.800 69.735 145.380 70.065 ;
        RECT 154.910 69.180 155.510 69.210 ;
        RECT 150.465 69.030 150.795 69.045 ;
        RECT 153.825 69.030 157.825 69.180 ;
        RECT 150.465 68.730 157.825 69.030 ;
        RECT 150.465 68.715 150.795 68.730 ;
        RECT 153.825 68.580 157.825 68.730 ;
        RECT 154.910 68.550 155.510 68.580 ;
        RECT 27.310 67.750 27.900 67.900 ;
        RECT 27.310 67.450 32.290 67.750 ;
        RECT 27.310 67.270 27.900 67.450 ;
        RECT 31.990 66.105 32.290 67.450 ;
        RECT 101.215 67.015 102.795 67.345 ;
        RECT 116.510 67.015 118.090 67.345 ;
        RECT 131.805 67.015 133.385 67.345 ;
        RECT 147.100 67.015 148.680 67.345 ;
        RECT 3.565 65.800 34.850 66.105 ;
        RECT 1.000 62.600 2.500 64.120 ;
        RECT 27.550 63.225 28.240 63.780 ;
        RECT 28.685 59.095 29.310 59.605 ;
        RECT 28.690 59.090 29.305 59.095 ;
        RECT 23.180 56.600 23.630 57.180 ;
        RECT 23.060 48.560 25.760 50.500 ;
        RECT 0.995 35.135 2.505 36.290 ;
        RECT 1.000 23.170 2.510 25.490 ;
        RECT 31.990 20.885 32.290 65.800 ;
        RECT 34.545 65.275 34.850 65.800 ;
        RECT 34.540 65.080 34.850 65.275 ;
        RECT 34.430 64.585 34.980 65.080 ;
        RECT 34.455 64.580 34.835 64.585 ;
        RECT 97.915 64.295 99.495 64.625 ;
        RECT 113.210 64.295 114.790 64.625 ;
        RECT 128.505 64.295 130.085 64.625 ;
        RECT 143.800 64.295 145.380 64.625 ;
        RECT 53.130 61.095 54.030 61.775 ;
        RECT 101.215 61.575 102.795 61.905 ;
        RECT 116.510 61.575 118.090 61.905 ;
        RECT 131.805 61.575 133.385 61.905 ;
        RECT 147.100 61.575 148.680 61.905 ;
        RECT 33.990 59.080 34.890 59.725 ;
        RECT 97.915 58.855 99.495 59.185 ;
        RECT 113.210 58.855 114.790 59.185 ;
        RECT 128.505 58.855 130.085 59.185 ;
        RECT 143.800 58.855 145.380 59.185 ;
        RECT 55.390 56.715 56.290 57.505 ;
        RECT 101.215 56.135 102.795 56.465 ;
        RECT 116.510 56.135 118.090 56.465 ;
        RECT 131.805 56.135 133.385 56.465 ;
        RECT 147.100 56.135 148.680 56.465 ;
        RECT 97.915 53.415 99.495 53.745 ;
        RECT 113.210 53.415 114.790 53.745 ;
        RECT 128.505 53.415 130.085 53.745 ;
        RECT 143.800 53.415 145.380 53.745 ;
        RECT 101.215 50.695 102.795 51.025 ;
        RECT 116.510 50.695 118.090 51.025 ;
        RECT 131.805 50.695 133.385 51.025 ;
        RECT 147.100 50.695 148.680 51.025 ;
        RECT 150.465 48.630 150.795 48.645 ;
        RECT 153.825 48.630 157.825 48.780 ;
        RECT 150.465 48.330 157.825 48.630 ;
        RECT 150.465 48.315 150.795 48.330 ;
        RECT 97.915 47.975 99.495 48.305 ;
        RECT 113.210 47.975 114.790 48.305 ;
        RECT 128.505 47.975 130.085 48.305 ;
        RECT 143.800 47.975 145.380 48.305 ;
        RECT 153.825 48.180 157.825 48.330 ;
        RECT 101.215 45.255 102.795 45.585 ;
        RECT 116.510 45.255 118.090 45.585 ;
        RECT 131.805 45.255 133.385 45.585 ;
        RECT 147.100 45.255 148.680 45.585 ;
        RECT 97.915 42.535 99.495 42.865 ;
        RECT 113.210 42.535 114.790 42.865 ;
        RECT 128.505 42.535 130.085 42.865 ;
        RECT 143.800 42.535 145.380 42.865 ;
        RECT 101.215 39.815 102.795 40.145 ;
        RECT 116.510 39.815 118.090 40.145 ;
        RECT 131.805 39.815 133.385 40.145 ;
        RECT 147.100 39.815 148.680 40.145 ;
        RECT 85.540 39.110 89.540 39.260 ;
        RECT 90.205 39.110 90.535 39.125 ;
        RECT 85.540 38.810 90.535 39.110 ;
        RECT 85.540 38.660 89.540 38.810 ;
        RECT 90.205 38.795 90.535 38.810 ;
        RECT 98.945 38.430 99.275 38.445 ;
        RECT 112.745 38.430 113.075 38.445 ;
        RECT 98.945 38.130 113.075 38.430 ;
        RECT 98.945 38.115 99.275 38.130 ;
        RECT 112.745 38.115 113.075 38.130 ;
        RECT 117.805 37.750 118.135 37.765 ;
        RECT 127.005 37.750 127.335 37.765 ;
        RECT 117.805 37.450 127.335 37.750 ;
        RECT 117.805 37.435 118.135 37.450 ;
        RECT 127.005 37.435 127.335 37.450 ;
        RECT 97.915 37.095 99.495 37.425 ;
        RECT 113.210 37.095 114.790 37.425 ;
        RECT 128.505 37.095 130.085 37.425 ;
        RECT 143.800 37.095 145.380 37.425 ;
        RECT 121.485 35.710 121.815 35.725 ;
        RECT 127.005 35.710 127.335 35.725 ;
        RECT 121.485 35.410 127.335 35.710 ;
        RECT 121.485 35.395 121.815 35.410 ;
        RECT 127.005 35.395 127.335 35.410 ;
        RECT 101.215 34.375 102.795 34.705 ;
        RECT 116.510 34.375 118.090 34.705 ;
        RECT 131.805 34.375 133.385 34.705 ;
        RECT 147.100 34.375 148.680 34.705 ;
        RECT 97.915 31.655 99.495 31.985 ;
        RECT 113.210 31.655 114.790 31.985 ;
        RECT 128.505 31.655 130.085 31.985 ;
        RECT 143.800 31.655 145.380 31.985 ;
        RECT 101.215 28.935 102.795 29.265 ;
        RECT 116.510 28.935 118.090 29.265 ;
        RECT 131.805 28.935 133.385 29.265 ;
        RECT 147.100 28.935 148.680 29.265 ;
        RECT 157.200 28.380 157.855 28.415 ;
        RECT 151.845 28.230 152.175 28.245 ;
        RECT 153.825 28.230 157.855 28.380 ;
        RECT 151.845 27.930 157.855 28.230 ;
        RECT 151.845 27.915 152.175 27.930 ;
        RECT 153.825 27.780 157.855 27.930 ;
        RECT 157.200 27.750 157.855 27.780 ;
        RECT 59.010 20.885 59.440 20.940 ;
        RECT 31.990 20.585 59.440 20.885 ;
        RECT 59.010 20.540 59.440 20.585 ;
        RECT 8.230 18.065 10.045 18.735 ;
        RECT 49.000 18.065 50.495 18.070 ;
        RECT 8.230 16.575 50.495 18.065 ;
        RECT 8.230 16.570 50.230 16.575 ;
        RECT 8.230 15.990 10.045 16.570 ;
        RECT 71.150 15.215 71.955 16.015 ;
        RECT 69.770 14.560 70.290 15.045 ;
        RECT 68.575 13.665 69.095 14.150 ;
        RECT 67.610 12.995 68.130 13.480 ;
        RECT 66.655 12.400 67.175 12.885 ;
        RECT 65.625 11.615 66.145 12.100 ;
        RECT 64.650 10.850 65.170 11.335 ;
        RECT 63.640 9.785 64.160 10.270 ;
        RECT 62.440 9.015 62.960 9.500 ;
        RECT 53.125 7.780 54.035 8.675 ;
        RECT 82.945 7.520 83.930 8.425 ;
        RECT 23.925 6.730 24.835 7.480 ;
        RECT 80.940 6.235 82.120 6.480 ;
        RECT 13.370 5.775 82.120 6.235 ;
        RECT 80.940 5.575 82.120 5.775 ;
      LAYER via3 ;
        RECT 154.780 223.130 155.350 223.815 ;
        RECT 84.910 222.545 85.260 222.895 ;
        RECT 88.580 222.550 88.930 222.900 ;
        RECT 66.565 220.495 66.885 220.815 ;
        RECT 70.205 220.535 70.525 220.855 ;
        RECT 147.325 220.850 147.975 221.450 ;
        RECT 46.555 218.905 46.875 219.225 ;
        RECT 44.575 217.615 44.895 217.935 ;
        RECT 143.635 218.935 144.285 219.585 ;
        RECT 139.955 216.755 140.605 217.405 ;
        RECT 153.630 216.785 154.220 217.375 ;
        RECT 136.295 215.090 136.945 215.740 ;
        RECT 153.870 215.120 154.460 215.710 ;
        RECT 4.200 213.295 4.520 213.630 ;
        RECT 62.905 213.320 63.225 213.640 ;
        RECT 1.470 194.160 2.020 194.710 ;
        RECT 1.365 82.730 2.055 83.240 ;
        RECT 157.230 220.830 157.820 221.420 ;
        RECT 155.985 218.965 156.575 219.555 ;
        RECT 35.255 153.405 35.575 155.525 ;
        RECT 20.380 149.800 20.730 150.150 ;
        RECT 35.255 149.805 35.575 151.925 ;
        RECT 24.120 145.940 26.240 146.260 ;
        RECT 35.255 146.205 35.575 148.325 ;
        RECT 25.545 143.440 26.260 144.195 ;
        RECT 21.045 142.955 21.395 143.305 ;
        RECT 35.255 142.605 35.575 144.725 ;
        RECT 35.255 139.005 35.575 141.125 ;
        RECT 35.255 135.405 35.575 137.525 ;
        RECT 35.255 131.805 35.575 133.925 ;
        RECT 35.255 128.205 35.575 130.325 ;
        RECT 35.255 124.605 35.575 126.725 ;
        RECT 76.525 194.270 76.845 194.590 ;
        RECT 76.925 194.270 77.245 194.590 ;
        RECT 77.325 194.270 77.645 194.590 ;
        RECT 77.725 194.270 78.045 194.590 ;
        RECT 88.600 194.270 88.920 194.590 ;
        RECT 89.000 194.270 89.320 194.590 ;
        RECT 89.400 194.270 89.720 194.590 ;
        RECT 89.800 194.270 90.120 194.590 ;
        RECT 100.675 194.270 100.995 194.590 ;
        RECT 101.075 194.270 101.395 194.590 ;
        RECT 101.475 194.270 101.795 194.590 ;
        RECT 101.875 194.270 102.195 194.590 ;
        RECT 112.750 194.270 113.070 194.590 ;
        RECT 113.150 194.270 113.470 194.590 ;
        RECT 113.550 194.270 113.870 194.590 ;
        RECT 113.950 194.270 114.270 194.590 ;
        RECT 79.825 191.550 80.145 191.870 ;
        RECT 80.225 191.550 80.545 191.870 ;
        RECT 80.625 191.550 80.945 191.870 ;
        RECT 81.025 191.550 81.345 191.870 ;
        RECT 91.900 191.550 92.220 191.870 ;
        RECT 92.300 191.550 92.620 191.870 ;
        RECT 92.700 191.550 93.020 191.870 ;
        RECT 93.100 191.550 93.420 191.870 ;
        RECT 103.975 191.550 104.295 191.870 ;
        RECT 104.375 191.550 104.695 191.870 ;
        RECT 104.775 191.550 105.095 191.870 ;
        RECT 105.175 191.550 105.495 191.870 ;
        RECT 116.050 191.550 116.370 191.870 ;
        RECT 116.450 191.550 116.770 191.870 ;
        RECT 116.850 191.550 117.170 191.870 ;
        RECT 117.250 191.550 117.570 191.870 ;
        RECT 67.325 189.035 67.645 189.355 ;
        RECT 76.525 188.830 76.845 189.150 ;
        RECT 76.925 188.830 77.245 189.150 ;
        RECT 77.325 188.830 77.645 189.150 ;
        RECT 77.725 188.830 78.045 189.150 ;
        RECT 88.600 188.830 88.920 189.150 ;
        RECT 89.000 188.830 89.320 189.150 ;
        RECT 89.400 188.830 89.720 189.150 ;
        RECT 89.800 188.830 90.120 189.150 ;
        RECT 100.675 188.830 100.995 189.150 ;
        RECT 101.075 188.830 101.395 189.150 ;
        RECT 101.475 188.830 101.795 189.150 ;
        RECT 101.875 188.830 102.195 189.150 ;
        RECT 112.750 188.830 113.070 189.150 ;
        RECT 113.150 188.830 113.470 189.150 ;
        RECT 113.550 188.830 113.870 189.150 ;
        RECT 113.950 188.830 114.270 189.150 ;
        RECT 128.945 189.030 129.545 189.630 ;
        RECT 79.825 186.110 80.145 186.430 ;
        RECT 80.225 186.110 80.545 186.430 ;
        RECT 80.625 186.110 80.945 186.430 ;
        RECT 81.025 186.110 81.345 186.430 ;
        RECT 91.900 186.110 92.220 186.430 ;
        RECT 92.300 186.110 92.620 186.430 ;
        RECT 92.700 186.110 93.020 186.430 ;
        RECT 93.100 186.110 93.420 186.430 ;
        RECT 103.975 186.110 104.295 186.430 ;
        RECT 104.375 186.110 104.695 186.430 ;
        RECT 104.775 186.110 105.095 186.430 ;
        RECT 105.175 186.110 105.495 186.430 ;
        RECT 116.050 186.110 116.370 186.430 ;
        RECT 116.450 186.110 116.770 186.430 ;
        RECT 116.850 186.110 117.170 186.430 ;
        RECT 117.250 186.110 117.570 186.430 ;
        RECT 76.525 183.390 76.845 183.710 ;
        RECT 76.925 183.390 77.245 183.710 ;
        RECT 77.325 183.390 77.645 183.710 ;
        RECT 77.725 183.390 78.045 183.710 ;
        RECT 88.600 183.390 88.920 183.710 ;
        RECT 89.000 183.390 89.320 183.710 ;
        RECT 89.400 183.390 89.720 183.710 ;
        RECT 89.800 183.390 90.120 183.710 ;
        RECT 100.675 183.390 100.995 183.710 ;
        RECT 101.075 183.390 101.395 183.710 ;
        RECT 101.475 183.390 101.795 183.710 ;
        RECT 101.875 183.390 102.195 183.710 ;
        RECT 112.750 183.390 113.070 183.710 ;
        RECT 113.150 183.390 113.470 183.710 ;
        RECT 113.550 183.390 113.870 183.710 ;
        RECT 113.950 183.390 114.270 183.710 ;
        RECT 79.825 180.670 80.145 180.990 ;
        RECT 80.225 180.670 80.545 180.990 ;
        RECT 80.625 180.670 80.945 180.990 ;
        RECT 81.025 180.670 81.345 180.990 ;
        RECT 91.900 180.670 92.220 180.990 ;
        RECT 92.300 180.670 92.620 180.990 ;
        RECT 92.700 180.670 93.020 180.990 ;
        RECT 93.100 180.670 93.420 180.990 ;
        RECT 103.975 180.670 104.295 180.990 ;
        RECT 104.375 180.670 104.695 180.990 ;
        RECT 104.775 180.670 105.095 180.990 ;
        RECT 105.175 180.670 105.495 180.990 ;
        RECT 116.050 180.670 116.370 180.990 ;
        RECT 116.450 180.670 116.770 180.990 ;
        RECT 116.850 180.670 117.170 180.990 ;
        RECT 117.250 180.670 117.570 180.990 ;
        RECT 76.525 177.950 76.845 178.270 ;
        RECT 76.925 177.950 77.245 178.270 ;
        RECT 77.325 177.950 77.645 178.270 ;
        RECT 77.725 177.950 78.045 178.270 ;
        RECT 88.600 177.950 88.920 178.270 ;
        RECT 89.000 177.950 89.320 178.270 ;
        RECT 89.400 177.950 89.720 178.270 ;
        RECT 89.800 177.950 90.120 178.270 ;
        RECT 100.675 177.950 100.995 178.270 ;
        RECT 101.075 177.950 101.395 178.270 ;
        RECT 101.475 177.950 101.795 178.270 ;
        RECT 101.875 177.950 102.195 178.270 ;
        RECT 112.750 177.950 113.070 178.270 ;
        RECT 113.150 177.950 113.470 178.270 ;
        RECT 113.550 177.950 113.870 178.270 ;
        RECT 113.950 177.950 114.270 178.270 ;
        RECT 79.825 175.230 80.145 175.550 ;
        RECT 80.225 175.230 80.545 175.550 ;
        RECT 80.625 175.230 80.945 175.550 ;
        RECT 81.025 175.230 81.345 175.550 ;
        RECT 91.900 175.230 92.220 175.550 ;
        RECT 92.300 175.230 92.620 175.550 ;
        RECT 92.700 175.230 93.020 175.550 ;
        RECT 93.100 175.230 93.420 175.550 ;
        RECT 103.975 175.230 104.295 175.550 ;
        RECT 104.375 175.230 104.695 175.550 ;
        RECT 104.775 175.230 105.095 175.550 ;
        RECT 105.175 175.230 105.495 175.550 ;
        RECT 116.050 175.230 116.370 175.550 ;
        RECT 116.450 175.230 116.770 175.550 ;
        RECT 116.850 175.230 117.170 175.550 ;
        RECT 117.250 175.230 117.570 175.550 ;
        RECT 76.525 172.510 76.845 172.830 ;
        RECT 76.925 172.510 77.245 172.830 ;
        RECT 77.325 172.510 77.645 172.830 ;
        RECT 77.725 172.510 78.045 172.830 ;
        RECT 88.600 172.510 88.920 172.830 ;
        RECT 89.000 172.510 89.320 172.830 ;
        RECT 89.400 172.510 89.720 172.830 ;
        RECT 89.800 172.510 90.120 172.830 ;
        RECT 100.675 172.510 100.995 172.830 ;
        RECT 101.075 172.510 101.395 172.830 ;
        RECT 101.475 172.510 101.795 172.830 ;
        RECT 101.875 172.510 102.195 172.830 ;
        RECT 112.750 172.510 113.070 172.830 ;
        RECT 113.150 172.510 113.470 172.830 ;
        RECT 113.550 172.510 113.870 172.830 ;
        RECT 113.950 172.510 114.270 172.830 ;
        RECT 79.825 169.790 80.145 170.110 ;
        RECT 80.225 169.790 80.545 170.110 ;
        RECT 80.625 169.790 80.945 170.110 ;
        RECT 81.025 169.790 81.345 170.110 ;
        RECT 91.900 169.790 92.220 170.110 ;
        RECT 92.300 169.790 92.620 170.110 ;
        RECT 92.700 169.790 93.020 170.110 ;
        RECT 93.100 169.790 93.420 170.110 ;
        RECT 103.975 169.790 104.295 170.110 ;
        RECT 104.375 169.790 104.695 170.110 ;
        RECT 104.775 169.790 105.095 170.110 ;
        RECT 105.175 169.790 105.495 170.110 ;
        RECT 116.050 169.790 116.370 170.110 ;
        RECT 116.450 169.790 116.770 170.110 ;
        RECT 116.850 169.790 117.170 170.110 ;
        RECT 117.250 169.790 117.570 170.110 ;
        RECT 76.525 167.070 76.845 167.390 ;
        RECT 76.925 167.070 77.245 167.390 ;
        RECT 77.325 167.070 77.645 167.390 ;
        RECT 77.725 167.070 78.045 167.390 ;
        RECT 88.600 167.070 88.920 167.390 ;
        RECT 89.000 167.070 89.320 167.390 ;
        RECT 89.400 167.070 89.720 167.390 ;
        RECT 89.800 167.070 90.120 167.390 ;
        RECT 100.675 167.070 100.995 167.390 ;
        RECT 101.075 167.070 101.395 167.390 ;
        RECT 101.475 167.070 101.795 167.390 ;
        RECT 101.875 167.070 102.195 167.390 ;
        RECT 112.750 167.070 113.070 167.390 ;
        RECT 113.150 167.070 113.470 167.390 ;
        RECT 113.550 167.070 113.870 167.390 ;
        RECT 113.950 167.070 114.270 167.390 ;
        RECT 79.825 164.350 80.145 164.670 ;
        RECT 80.225 164.350 80.545 164.670 ;
        RECT 80.625 164.350 80.945 164.670 ;
        RECT 81.025 164.350 81.345 164.670 ;
        RECT 91.900 164.350 92.220 164.670 ;
        RECT 92.300 164.350 92.620 164.670 ;
        RECT 92.700 164.350 93.020 164.670 ;
        RECT 93.100 164.350 93.420 164.670 ;
        RECT 103.975 164.350 104.295 164.670 ;
        RECT 104.375 164.350 104.695 164.670 ;
        RECT 104.775 164.350 105.095 164.670 ;
        RECT 105.175 164.350 105.495 164.670 ;
        RECT 116.050 164.350 116.370 164.670 ;
        RECT 116.450 164.350 116.770 164.670 ;
        RECT 116.850 164.350 117.170 164.670 ;
        RECT 117.250 164.350 117.570 164.670 ;
        RECT 76.525 161.630 76.845 161.950 ;
        RECT 76.925 161.630 77.245 161.950 ;
        RECT 77.325 161.630 77.645 161.950 ;
        RECT 77.725 161.630 78.045 161.950 ;
        RECT 88.600 161.630 88.920 161.950 ;
        RECT 89.000 161.630 89.320 161.950 ;
        RECT 89.400 161.630 89.720 161.950 ;
        RECT 89.800 161.630 90.120 161.950 ;
        RECT 100.675 161.630 100.995 161.950 ;
        RECT 101.075 161.630 101.395 161.950 ;
        RECT 101.475 161.630 101.795 161.950 ;
        RECT 101.875 161.630 102.195 161.950 ;
        RECT 112.750 161.630 113.070 161.950 ;
        RECT 113.150 161.630 113.470 161.950 ;
        RECT 113.550 161.630 113.870 161.950 ;
        RECT 113.950 161.630 114.270 161.950 ;
        RECT 79.825 158.910 80.145 159.230 ;
        RECT 80.225 158.910 80.545 159.230 ;
        RECT 80.625 158.910 80.945 159.230 ;
        RECT 81.025 158.910 81.345 159.230 ;
        RECT 91.900 158.910 92.220 159.230 ;
        RECT 92.300 158.910 92.620 159.230 ;
        RECT 92.700 158.910 93.020 159.230 ;
        RECT 93.100 158.910 93.420 159.230 ;
        RECT 103.975 158.910 104.295 159.230 ;
        RECT 104.375 158.910 104.695 159.230 ;
        RECT 104.775 158.910 105.095 159.230 ;
        RECT 105.175 158.910 105.495 159.230 ;
        RECT 116.050 158.910 116.370 159.230 ;
        RECT 116.450 158.910 116.770 159.230 ;
        RECT 116.850 158.910 117.170 159.230 ;
        RECT 117.250 158.910 117.570 159.230 ;
        RECT 76.525 156.190 76.845 156.510 ;
        RECT 76.925 156.190 77.245 156.510 ;
        RECT 77.325 156.190 77.645 156.510 ;
        RECT 77.725 156.190 78.045 156.510 ;
        RECT 88.600 156.190 88.920 156.510 ;
        RECT 89.000 156.190 89.320 156.510 ;
        RECT 89.400 156.190 89.720 156.510 ;
        RECT 89.800 156.190 90.120 156.510 ;
        RECT 100.675 156.190 100.995 156.510 ;
        RECT 101.075 156.190 101.395 156.510 ;
        RECT 101.475 156.190 101.795 156.510 ;
        RECT 101.875 156.190 102.195 156.510 ;
        RECT 112.750 156.190 113.070 156.510 ;
        RECT 113.150 156.190 113.470 156.510 ;
        RECT 113.550 156.190 113.870 156.510 ;
        RECT 113.950 156.190 114.270 156.510 ;
        RECT 49.390 147.925 49.920 148.455 ;
        RECT 79.825 153.470 80.145 153.790 ;
        RECT 80.225 153.470 80.545 153.790 ;
        RECT 80.625 153.470 80.945 153.790 ;
        RECT 81.025 153.470 81.345 153.790 ;
        RECT 91.900 153.470 92.220 153.790 ;
        RECT 92.300 153.470 92.620 153.790 ;
        RECT 92.700 153.470 93.020 153.790 ;
        RECT 93.100 153.470 93.420 153.790 ;
        RECT 103.975 153.470 104.295 153.790 ;
        RECT 104.375 153.470 104.695 153.790 ;
        RECT 104.775 153.470 105.095 153.790 ;
        RECT 105.175 153.470 105.495 153.790 ;
        RECT 116.050 153.470 116.370 153.790 ;
        RECT 116.450 153.470 116.770 153.790 ;
        RECT 116.850 153.470 117.170 153.790 ;
        RECT 117.250 153.470 117.570 153.790 ;
        RECT 132.540 153.670 133.140 154.270 ;
        RECT 76.525 150.750 76.845 151.070 ;
        RECT 76.925 150.750 77.245 151.070 ;
        RECT 77.325 150.750 77.645 151.070 ;
        RECT 77.725 150.750 78.045 151.070 ;
        RECT 88.600 150.750 88.920 151.070 ;
        RECT 89.000 150.750 89.320 151.070 ;
        RECT 89.400 150.750 89.720 151.070 ;
        RECT 89.800 150.750 90.120 151.070 ;
        RECT 100.675 150.750 100.995 151.070 ;
        RECT 101.075 150.750 101.395 151.070 ;
        RECT 101.475 150.750 101.795 151.070 ;
        RECT 101.875 150.750 102.195 151.070 ;
        RECT 112.750 150.750 113.070 151.070 ;
        RECT 113.150 150.750 113.470 151.070 ;
        RECT 113.550 150.750 113.870 151.070 ;
        RECT 113.950 150.750 114.270 151.070 ;
        RECT 79.825 148.030 80.145 148.350 ;
        RECT 80.225 148.030 80.545 148.350 ;
        RECT 80.625 148.030 80.945 148.350 ;
        RECT 81.025 148.030 81.345 148.350 ;
        RECT 91.900 148.030 92.220 148.350 ;
        RECT 92.300 148.030 92.620 148.350 ;
        RECT 92.700 148.030 93.020 148.350 ;
        RECT 93.100 148.030 93.420 148.350 ;
        RECT 103.975 148.030 104.295 148.350 ;
        RECT 104.375 148.030 104.695 148.350 ;
        RECT 104.775 148.030 105.095 148.350 ;
        RECT 105.175 148.030 105.495 148.350 ;
        RECT 116.050 148.030 116.370 148.350 ;
        RECT 116.450 148.030 116.770 148.350 ;
        RECT 116.850 148.030 117.170 148.350 ;
        RECT 117.250 148.030 117.570 148.350 ;
        RECT 80.280 139.075 81.170 139.965 ;
        RECT 110.375 139.260 110.885 139.820 ;
        RECT 79.015 124.505 79.975 125.315 ;
        RECT 35.035 115.435 35.355 117.555 ;
        RECT 20.160 111.830 20.510 112.180 ;
        RECT 35.035 111.835 35.355 113.955 ;
        RECT 23.900 107.970 26.020 108.290 ;
        RECT 35.035 108.235 35.355 110.355 ;
        RECT 25.325 105.470 26.040 106.225 ;
        RECT 20.825 104.985 21.175 105.335 ;
        RECT 35.035 104.635 35.355 106.755 ;
        RECT 35.035 101.035 35.355 103.155 ;
        RECT 35.035 97.435 35.355 99.555 ;
        RECT 35.035 93.835 35.355 95.955 ;
        RECT 35.035 90.235 35.355 92.355 ;
        RECT 35.035 86.635 35.355 88.755 ;
        RECT 46.540 121.885 46.890 122.235 ;
        RECT 44.560 88.945 44.910 89.295 ;
        RECT 49.350 88.610 50.010 89.310 ;
        RECT 152.035 135.275 152.685 135.875 ;
        RECT 101.245 88.780 101.565 89.100 ;
        RECT 101.645 88.780 101.965 89.100 ;
        RECT 102.045 88.780 102.365 89.100 ;
        RECT 102.445 88.780 102.765 89.100 ;
        RECT 116.540 88.780 116.860 89.100 ;
        RECT 116.940 88.780 117.260 89.100 ;
        RECT 117.340 88.780 117.660 89.100 ;
        RECT 117.740 88.780 118.060 89.100 ;
        RECT 131.835 88.780 132.155 89.100 ;
        RECT 132.235 88.780 132.555 89.100 ;
        RECT 132.635 88.780 132.955 89.100 ;
        RECT 133.035 88.780 133.355 89.100 ;
        RECT 147.130 88.780 147.450 89.100 ;
        RECT 147.530 88.780 147.850 89.100 ;
        RECT 147.930 88.780 148.250 89.100 ;
        RECT 148.330 88.780 148.650 89.100 ;
        RECT 153.865 88.980 154.465 89.580 ;
        RECT 97.945 86.060 98.265 86.380 ;
        RECT 98.345 86.060 98.665 86.380 ;
        RECT 98.745 86.060 99.065 86.380 ;
        RECT 99.145 86.060 99.465 86.380 ;
        RECT 113.240 86.060 113.560 86.380 ;
        RECT 113.640 86.060 113.960 86.380 ;
        RECT 114.040 86.060 114.360 86.380 ;
        RECT 114.440 86.060 114.760 86.380 ;
        RECT 128.535 86.060 128.855 86.380 ;
        RECT 128.935 86.060 129.255 86.380 ;
        RECT 129.335 86.060 129.655 86.380 ;
        RECT 129.735 86.060 130.055 86.380 ;
        RECT 143.830 86.060 144.150 86.380 ;
        RECT 144.230 86.060 144.550 86.380 ;
        RECT 144.630 86.060 144.950 86.380 ;
        RECT 145.030 86.060 145.350 86.380 ;
        RECT 101.245 83.340 101.565 83.660 ;
        RECT 101.645 83.340 101.965 83.660 ;
        RECT 102.045 83.340 102.365 83.660 ;
        RECT 102.445 83.340 102.765 83.660 ;
        RECT 116.540 83.340 116.860 83.660 ;
        RECT 116.940 83.340 117.260 83.660 ;
        RECT 117.340 83.340 117.660 83.660 ;
        RECT 117.740 83.340 118.060 83.660 ;
        RECT 131.835 83.340 132.155 83.660 ;
        RECT 132.235 83.340 132.555 83.660 ;
        RECT 132.635 83.340 132.955 83.660 ;
        RECT 133.035 83.340 133.355 83.660 ;
        RECT 147.130 83.340 147.450 83.660 ;
        RECT 147.530 83.340 147.850 83.660 ;
        RECT 147.930 83.340 148.250 83.660 ;
        RECT 148.330 83.340 148.650 83.660 ;
        RECT 97.945 80.620 98.265 80.940 ;
        RECT 98.345 80.620 98.665 80.940 ;
        RECT 98.745 80.620 99.065 80.940 ;
        RECT 99.145 80.620 99.465 80.940 ;
        RECT 113.240 80.620 113.560 80.940 ;
        RECT 113.640 80.620 113.960 80.940 ;
        RECT 114.040 80.620 114.360 80.940 ;
        RECT 114.440 80.620 114.760 80.940 ;
        RECT 128.535 80.620 128.855 80.940 ;
        RECT 128.935 80.620 129.255 80.940 ;
        RECT 129.335 80.620 129.655 80.940 ;
        RECT 129.735 80.620 130.055 80.940 ;
        RECT 143.830 80.620 144.150 80.940 ;
        RECT 144.230 80.620 144.550 80.940 ;
        RECT 144.630 80.620 144.950 80.940 ;
        RECT 145.030 80.620 145.350 80.940 ;
        RECT 101.245 77.900 101.565 78.220 ;
        RECT 101.645 77.900 101.965 78.220 ;
        RECT 102.045 77.900 102.365 78.220 ;
        RECT 102.445 77.900 102.765 78.220 ;
        RECT 116.540 77.900 116.860 78.220 ;
        RECT 116.940 77.900 117.260 78.220 ;
        RECT 117.340 77.900 117.660 78.220 ;
        RECT 117.740 77.900 118.060 78.220 ;
        RECT 131.835 77.900 132.155 78.220 ;
        RECT 132.235 77.900 132.555 78.220 ;
        RECT 132.635 77.900 132.955 78.220 ;
        RECT 133.035 77.900 133.355 78.220 ;
        RECT 147.130 77.900 147.450 78.220 ;
        RECT 147.530 77.900 147.850 78.220 ;
        RECT 147.930 77.900 148.250 78.220 ;
        RECT 148.330 77.900 148.650 78.220 ;
        RECT 97.945 75.180 98.265 75.500 ;
        RECT 98.345 75.180 98.665 75.500 ;
        RECT 98.745 75.180 99.065 75.500 ;
        RECT 99.145 75.180 99.465 75.500 ;
        RECT 113.240 75.180 113.560 75.500 ;
        RECT 113.640 75.180 113.960 75.500 ;
        RECT 114.040 75.180 114.360 75.500 ;
        RECT 114.440 75.180 114.760 75.500 ;
        RECT 128.535 75.180 128.855 75.500 ;
        RECT 128.935 75.180 129.255 75.500 ;
        RECT 129.335 75.180 129.655 75.500 ;
        RECT 129.735 75.180 130.055 75.500 ;
        RECT 143.830 75.180 144.150 75.500 ;
        RECT 144.230 75.180 144.550 75.500 ;
        RECT 144.630 75.180 144.950 75.500 ;
        RECT 145.030 75.180 145.350 75.500 ;
        RECT 101.245 72.460 101.565 72.780 ;
        RECT 101.645 72.460 101.965 72.780 ;
        RECT 102.045 72.460 102.365 72.780 ;
        RECT 102.445 72.460 102.765 72.780 ;
        RECT 116.540 72.460 116.860 72.780 ;
        RECT 116.940 72.460 117.260 72.780 ;
        RECT 117.340 72.460 117.660 72.780 ;
        RECT 117.740 72.460 118.060 72.780 ;
        RECT 131.835 72.460 132.155 72.780 ;
        RECT 132.235 72.460 132.555 72.780 ;
        RECT 132.635 72.460 132.955 72.780 ;
        RECT 133.035 72.460 133.355 72.780 ;
        RECT 147.130 72.460 147.450 72.780 ;
        RECT 147.530 72.460 147.850 72.780 ;
        RECT 147.930 72.460 148.250 72.780 ;
        RECT 148.330 72.460 148.650 72.780 ;
        RECT 27.570 69.705 27.905 70.030 ;
        RECT 97.945 69.740 98.265 70.060 ;
        RECT 98.345 69.740 98.665 70.060 ;
        RECT 98.745 69.740 99.065 70.060 ;
        RECT 99.145 69.740 99.465 70.060 ;
        RECT 113.240 69.740 113.560 70.060 ;
        RECT 113.640 69.740 113.960 70.060 ;
        RECT 114.040 69.740 114.360 70.060 ;
        RECT 114.440 69.740 114.760 70.060 ;
        RECT 128.535 69.740 128.855 70.060 ;
        RECT 128.935 69.740 129.255 70.060 ;
        RECT 129.335 69.740 129.655 70.060 ;
        RECT 129.735 69.740 130.055 70.060 ;
        RECT 143.830 69.740 144.150 70.060 ;
        RECT 144.230 69.740 144.550 70.060 ;
        RECT 144.630 69.740 144.950 70.060 ;
        RECT 145.030 69.740 145.350 70.060 ;
        RECT 49.470 68.890 50.090 69.680 ;
        RECT 154.910 68.580 155.510 69.180 ;
        RECT 101.245 67.020 101.565 67.340 ;
        RECT 101.645 67.020 101.965 67.340 ;
        RECT 102.045 67.020 102.365 67.340 ;
        RECT 102.445 67.020 102.765 67.340 ;
        RECT 116.540 67.020 116.860 67.340 ;
        RECT 116.940 67.020 117.260 67.340 ;
        RECT 117.340 67.020 117.660 67.340 ;
        RECT 117.740 67.020 118.060 67.340 ;
        RECT 131.835 67.020 132.155 67.340 ;
        RECT 132.235 67.020 132.555 67.340 ;
        RECT 132.635 67.020 132.955 67.340 ;
        RECT 133.035 67.020 133.355 67.340 ;
        RECT 147.130 67.020 147.450 67.340 ;
        RECT 147.530 67.020 147.850 67.340 ;
        RECT 147.930 67.020 148.250 67.340 ;
        RECT 148.330 67.020 148.650 67.340 ;
        RECT 1.320 62.900 1.940 63.690 ;
        RECT 27.730 63.340 28.065 63.665 ;
        RECT 28.780 59.195 29.190 59.545 ;
        RECT 23.630 48.930 25.220 50.170 ;
        RECT 1.280 35.295 2.220 36.155 ;
        RECT 1.280 23.810 2.220 24.670 ;
        RECT 97.945 64.300 98.265 64.620 ;
        RECT 98.345 64.300 98.665 64.620 ;
        RECT 98.745 64.300 99.065 64.620 ;
        RECT 99.145 64.300 99.465 64.620 ;
        RECT 113.240 64.300 113.560 64.620 ;
        RECT 113.640 64.300 113.960 64.620 ;
        RECT 114.040 64.300 114.360 64.620 ;
        RECT 114.440 64.300 114.760 64.620 ;
        RECT 128.535 64.300 128.855 64.620 ;
        RECT 128.935 64.300 129.255 64.620 ;
        RECT 129.335 64.300 129.655 64.620 ;
        RECT 129.735 64.300 130.055 64.620 ;
        RECT 143.830 64.300 144.150 64.620 ;
        RECT 144.230 64.300 144.550 64.620 ;
        RECT 144.630 64.300 144.950 64.620 ;
        RECT 145.030 64.300 145.350 64.620 ;
        RECT 53.395 61.225 53.760 61.605 ;
        RECT 101.245 61.580 101.565 61.900 ;
        RECT 101.645 61.580 101.965 61.900 ;
        RECT 102.045 61.580 102.365 61.900 ;
        RECT 102.445 61.580 102.765 61.900 ;
        RECT 116.540 61.580 116.860 61.900 ;
        RECT 116.940 61.580 117.260 61.900 ;
        RECT 117.340 61.580 117.660 61.900 ;
        RECT 117.740 61.580 118.060 61.900 ;
        RECT 131.835 61.580 132.155 61.900 ;
        RECT 132.235 61.580 132.555 61.900 ;
        RECT 132.635 61.580 132.955 61.900 ;
        RECT 133.035 61.580 133.355 61.900 ;
        RECT 147.130 61.580 147.450 61.900 ;
        RECT 147.530 61.580 147.850 61.900 ;
        RECT 147.930 61.580 148.250 61.900 ;
        RECT 148.330 61.580 148.650 61.900 ;
        RECT 34.220 59.225 34.670 59.575 ;
        RECT 97.945 58.860 98.265 59.180 ;
        RECT 98.345 58.860 98.665 59.180 ;
        RECT 98.745 58.860 99.065 59.180 ;
        RECT 99.145 58.860 99.465 59.180 ;
        RECT 113.240 58.860 113.560 59.180 ;
        RECT 113.640 58.860 113.960 59.180 ;
        RECT 114.040 58.860 114.360 59.180 ;
        RECT 114.440 58.860 114.760 59.180 ;
        RECT 128.535 58.860 128.855 59.180 ;
        RECT 128.935 58.860 129.255 59.180 ;
        RECT 129.335 58.860 129.655 59.180 ;
        RECT 129.735 58.860 130.055 59.180 ;
        RECT 143.830 58.860 144.150 59.180 ;
        RECT 144.230 58.860 144.550 59.180 ;
        RECT 144.630 58.860 144.950 59.180 ;
        RECT 145.030 58.860 145.350 59.180 ;
        RECT 55.655 56.860 56.090 57.345 ;
        RECT 101.245 56.140 101.565 56.460 ;
        RECT 101.645 56.140 101.965 56.460 ;
        RECT 102.045 56.140 102.365 56.460 ;
        RECT 102.445 56.140 102.765 56.460 ;
        RECT 116.540 56.140 116.860 56.460 ;
        RECT 116.940 56.140 117.260 56.460 ;
        RECT 117.340 56.140 117.660 56.460 ;
        RECT 117.740 56.140 118.060 56.460 ;
        RECT 131.835 56.140 132.155 56.460 ;
        RECT 132.235 56.140 132.555 56.460 ;
        RECT 132.635 56.140 132.955 56.460 ;
        RECT 133.035 56.140 133.355 56.460 ;
        RECT 147.130 56.140 147.450 56.460 ;
        RECT 147.530 56.140 147.850 56.460 ;
        RECT 147.930 56.140 148.250 56.460 ;
        RECT 148.330 56.140 148.650 56.460 ;
        RECT 97.945 53.420 98.265 53.740 ;
        RECT 98.345 53.420 98.665 53.740 ;
        RECT 98.745 53.420 99.065 53.740 ;
        RECT 99.145 53.420 99.465 53.740 ;
        RECT 113.240 53.420 113.560 53.740 ;
        RECT 113.640 53.420 113.960 53.740 ;
        RECT 114.040 53.420 114.360 53.740 ;
        RECT 114.440 53.420 114.760 53.740 ;
        RECT 128.535 53.420 128.855 53.740 ;
        RECT 128.935 53.420 129.255 53.740 ;
        RECT 129.335 53.420 129.655 53.740 ;
        RECT 129.735 53.420 130.055 53.740 ;
        RECT 143.830 53.420 144.150 53.740 ;
        RECT 144.230 53.420 144.550 53.740 ;
        RECT 144.630 53.420 144.950 53.740 ;
        RECT 145.030 53.420 145.350 53.740 ;
        RECT 101.245 50.700 101.565 51.020 ;
        RECT 101.645 50.700 101.965 51.020 ;
        RECT 102.045 50.700 102.365 51.020 ;
        RECT 102.445 50.700 102.765 51.020 ;
        RECT 116.540 50.700 116.860 51.020 ;
        RECT 116.940 50.700 117.260 51.020 ;
        RECT 117.340 50.700 117.660 51.020 ;
        RECT 117.740 50.700 118.060 51.020 ;
        RECT 131.835 50.700 132.155 51.020 ;
        RECT 132.235 50.700 132.555 51.020 ;
        RECT 132.635 50.700 132.955 51.020 ;
        RECT 133.035 50.700 133.355 51.020 ;
        RECT 147.130 50.700 147.450 51.020 ;
        RECT 147.530 50.700 147.850 51.020 ;
        RECT 147.930 50.700 148.250 51.020 ;
        RECT 148.330 50.700 148.650 51.020 ;
        RECT 97.945 47.980 98.265 48.300 ;
        RECT 98.345 47.980 98.665 48.300 ;
        RECT 98.745 47.980 99.065 48.300 ;
        RECT 99.145 47.980 99.465 48.300 ;
        RECT 113.240 47.980 113.560 48.300 ;
        RECT 113.640 47.980 113.960 48.300 ;
        RECT 114.040 47.980 114.360 48.300 ;
        RECT 114.440 47.980 114.760 48.300 ;
        RECT 128.535 47.980 128.855 48.300 ;
        RECT 128.935 47.980 129.255 48.300 ;
        RECT 129.335 47.980 129.655 48.300 ;
        RECT 129.735 47.980 130.055 48.300 ;
        RECT 143.830 47.980 144.150 48.300 ;
        RECT 144.230 47.980 144.550 48.300 ;
        RECT 144.630 47.980 144.950 48.300 ;
        RECT 145.030 47.980 145.350 48.300 ;
        RECT 155.980 48.180 156.580 48.780 ;
        RECT 101.245 45.260 101.565 45.580 ;
        RECT 101.645 45.260 101.965 45.580 ;
        RECT 102.045 45.260 102.365 45.580 ;
        RECT 102.445 45.260 102.765 45.580 ;
        RECT 116.540 45.260 116.860 45.580 ;
        RECT 116.940 45.260 117.260 45.580 ;
        RECT 117.340 45.260 117.660 45.580 ;
        RECT 117.740 45.260 118.060 45.580 ;
        RECT 131.835 45.260 132.155 45.580 ;
        RECT 132.235 45.260 132.555 45.580 ;
        RECT 132.635 45.260 132.955 45.580 ;
        RECT 133.035 45.260 133.355 45.580 ;
        RECT 147.130 45.260 147.450 45.580 ;
        RECT 147.530 45.260 147.850 45.580 ;
        RECT 147.930 45.260 148.250 45.580 ;
        RECT 148.330 45.260 148.650 45.580 ;
        RECT 97.945 42.540 98.265 42.860 ;
        RECT 98.345 42.540 98.665 42.860 ;
        RECT 98.745 42.540 99.065 42.860 ;
        RECT 99.145 42.540 99.465 42.860 ;
        RECT 113.240 42.540 113.560 42.860 ;
        RECT 113.640 42.540 113.960 42.860 ;
        RECT 114.040 42.540 114.360 42.860 ;
        RECT 114.440 42.540 114.760 42.860 ;
        RECT 128.535 42.540 128.855 42.860 ;
        RECT 128.935 42.540 129.255 42.860 ;
        RECT 129.335 42.540 129.655 42.860 ;
        RECT 129.735 42.540 130.055 42.860 ;
        RECT 143.830 42.540 144.150 42.860 ;
        RECT 144.230 42.540 144.550 42.860 ;
        RECT 144.630 42.540 144.950 42.860 ;
        RECT 145.030 42.540 145.350 42.860 ;
        RECT 101.245 39.820 101.565 40.140 ;
        RECT 101.645 39.820 101.965 40.140 ;
        RECT 102.045 39.820 102.365 40.140 ;
        RECT 102.445 39.820 102.765 40.140 ;
        RECT 116.540 39.820 116.860 40.140 ;
        RECT 116.940 39.820 117.260 40.140 ;
        RECT 117.340 39.820 117.660 40.140 ;
        RECT 117.740 39.820 118.060 40.140 ;
        RECT 131.835 39.820 132.155 40.140 ;
        RECT 132.235 39.820 132.555 40.140 ;
        RECT 132.635 39.820 132.955 40.140 ;
        RECT 133.035 39.820 133.355 40.140 ;
        RECT 147.130 39.820 147.450 40.140 ;
        RECT 147.530 39.820 147.850 40.140 ;
        RECT 147.930 39.820 148.250 40.140 ;
        RECT 148.330 39.820 148.650 40.140 ;
        RECT 97.945 37.100 98.265 37.420 ;
        RECT 98.345 37.100 98.665 37.420 ;
        RECT 98.745 37.100 99.065 37.420 ;
        RECT 99.145 37.100 99.465 37.420 ;
        RECT 113.240 37.100 113.560 37.420 ;
        RECT 113.640 37.100 113.960 37.420 ;
        RECT 114.040 37.100 114.360 37.420 ;
        RECT 114.440 37.100 114.760 37.420 ;
        RECT 128.535 37.100 128.855 37.420 ;
        RECT 128.935 37.100 129.255 37.420 ;
        RECT 129.335 37.100 129.655 37.420 ;
        RECT 129.735 37.100 130.055 37.420 ;
        RECT 143.830 37.100 144.150 37.420 ;
        RECT 144.230 37.100 144.550 37.420 ;
        RECT 144.630 37.100 144.950 37.420 ;
        RECT 145.030 37.100 145.350 37.420 ;
        RECT 101.245 34.380 101.565 34.700 ;
        RECT 101.645 34.380 101.965 34.700 ;
        RECT 102.045 34.380 102.365 34.700 ;
        RECT 102.445 34.380 102.765 34.700 ;
        RECT 116.540 34.380 116.860 34.700 ;
        RECT 116.940 34.380 117.260 34.700 ;
        RECT 117.340 34.380 117.660 34.700 ;
        RECT 117.740 34.380 118.060 34.700 ;
        RECT 131.835 34.380 132.155 34.700 ;
        RECT 132.235 34.380 132.555 34.700 ;
        RECT 132.635 34.380 132.955 34.700 ;
        RECT 133.035 34.380 133.355 34.700 ;
        RECT 147.130 34.380 147.450 34.700 ;
        RECT 147.530 34.380 147.850 34.700 ;
        RECT 147.930 34.380 148.250 34.700 ;
        RECT 148.330 34.380 148.650 34.700 ;
        RECT 97.945 31.660 98.265 31.980 ;
        RECT 98.345 31.660 98.665 31.980 ;
        RECT 98.745 31.660 99.065 31.980 ;
        RECT 99.145 31.660 99.465 31.980 ;
        RECT 113.240 31.660 113.560 31.980 ;
        RECT 113.640 31.660 113.960 31.980 ;
        RECT 114.040 31.660 114.360 31.980 ;
        RECT 114.440 31.660 114.760 31.980 ;
        RECT 128.535 31.660 128.855 31.980 ;
        RECT 128.935 31.660 129.255 31.980 ;
        RECT 129.335 31.660 129.655 31.980 ;
        RECT 129.735 31.660 130.055 31.980 ;
        RECT 143.830 31.660 144.150 31.980 ;
        RECT 144.230 31.660 144.550 31.980 ;
        RECT 144.630 31.660 144.950 31.980 ;
        RECT 145.030 31.660 145.350 31.980 ;
        RECT 101.245 28.940 101.565 29.260 ;
        RECT 101.645 28.940 101.965 29.260 ;
        RECT 102.045 28.940 102.365 29.260 ;
        RECT 102.445 28.940 102.765 29.260 ;
        RECT 116.540 28.940 116.860 29.260 ;
        RECT 116.940 28.940 117.260 29.260 ;
        RECT 117.340 28.940 117.660 29.260 ;
        RECT 117.740 28.940 118.060 29.260 ;
        RECT 131.835 28.940 132.155 29.260 ;
        RECT 132.235 28.940 132.555 29.260 ;
        RECT 132.635 28.940 132.955 29.260 ;
        RECT 133.035 28.940 133.355 29.260 ;
        RECT 147.130 28.940 147.450 29.260 ;
        RECT 147.530 28.940 147.850 29.260 ;
        RECT 147.930 28.940 148.250 29.260 ;
        RECT 148.330 28.940 148.650 29.260 ;
        RECT 157.225 27.780 157.825 28.380 ;
        RECT 49.375 16.815 50.220 17.730 ;
        RECT 71.320 15.340 71.670 15.690 ;
        RECT 69.860 14.635 70.210 14.985 ;
        RECT 68.655 13.725 69.005 14.075 ;
        RECT 67.700 13.065 68.050 13.415 ;
        RECT 66.745 12.475 67.095 12.825 ;
        RECT 65.720 11.675 66.070 12.025 ;
        RECT 64.735 10.930 65.085 11.280 ;
        RECT 63.735 9.855 64.085 10.205 ;
        RECT 62.515 9.085 62.865 9.435 ;
        RECT 53.335 8.005 53.805 8.460 ;
        RECT 83.210 7.760 83.645 8.180 ;
        RECT 24.180 6.915 24.550 7.270 ;
        RECT 13.685 5.885 14.005 6.210 ;
        RECT 81.240 5.755 81.730 6.215 ;
      LAYER met4 ;
        RECT 66.850 224.760 66.875 225.050 ;
        RECT 33.430 224.440 33.730 224.760 ;
        RECT 46.550 218.900 46.880 219.230 ;
        RECT 44.570 217.610 44.900 217.940 ;
        RECT 4.105 213.265 4.550 213.665 ;
        RECT 2.500 193.685 2.505 195.185 ;
        RECT 4.210 59.465 4.520 213.265 ;
        RECT 9.125 157.330 33.275 157.850 ;
        RECT 9.125 74.220 9.645 157.330 ;
        RECT 32.755 156.435 33.275 157.330 ;
        RECT 32.750 156.125 33.275 156.435 ;
        RECT 32.755 155.270 33.275 156.125 ;
        RECT 32.210 154.670 33.820 155.270 ;
        RECT 28.915 154.030 33.820 154.670 ;
        RECT 20.375 149.795 20.735 150.155 ;
        RECT 20.405 148.995 20.720 149.795 ;
        RECT 24.375 148.995 25.985 149.305 ;
        RECT 20.340 148.475 25.985 148.995 ;
        RECT 20.350 148.470 25.985 148.475 ;
        RECT 20.350 143.280 20.650 148.470 ;
        RECT 24.375 147.695 25.985 148.470 ;
        RECT 24.040 145.860 26.320 146.340 ;
        RECT 25.335 144.155 26.440 144.355 ;
        RECT 28.915 144.155 29.555 154.030 ;
        RECT 32.210 153.660 33.820 154.030 ;
        RECT 32.755 151.670 33.275 153.660 ;
        RECT 32.210 150.060 33.820 151.670 ;
        RECT 32.755 148.070 33.275 150.060 ;
        RECT 32.210 146.460 33.820 148.070 ;
        RECT 32.755 144.470 33.275 146.460 ;
        RECT 25.335 143.515 29.555 144.155 ;
        RECT 21.040 143.280 21.400 143.310 ;
        RECT 20.350 142.980 21.400 143.280 ;
        RECT 25.335 143.245 26.440 143.515 ;
        RECT 21.040 142.950 21.400 142.980 ;
        RECT 32.210 142.860 33.820 144.470 ;
        RECT 32.755 140.870 33.275 142.860 ;
        RECT 32.210 139.260 33.820 140.870 ;
        RECT 32.755 137.270 33.275 139.260 ;
        RECT 32.210 135.660 33.820 137.270 ;
        RECT 32.755 133.670 33.275 135.660 ;
        RECT 32.210 132.060 33.820 133.670 ;
        RECT 32.755 130.070 33.275 132.060 ;
        RECT 32.210 128.460 33.820 130.070 ;
        RECT 32.755 126.470 33.275 128.460 ;
        RECT 32.210 124.860 33.820 126.470 ;
        RECT 32.755 123.865 33.275 124.860 ;
        RECT 35.155 123.865 35.675 156.265 ;
        RECT 32.535 120.420 39.110 120.940 ;
        RECT 32.535 117.300 33.055 120.420 ;
        RECT 31.990 116.700 33.600 117.300 ;
        RECT 28.695 116.060 33.600 116.700 ;
        RECT 20.155 111.825 20.515 112.185 ;
        RECT 20.185 111.025 20.500 111.825 ;
        RECT 24.155 111.025 25.765 111.335 ;
        RECT 20.120 110.505 25.765 111.025 ;
        RECT 20.130 110.500 25.765 110.505 ;
        RECT 20.130 105.310 20.430 110.500 ;
        RECT 24.155 109.725 25.765 110.500 ;
        RECT 23.820 107.890 26.100 108.370 ;
        RECT 25.115 106.185 26.220 106.385 ;
        RECT 28.695 106.185 29.335 116.060 ;
        RECT 31.990 115.690 33.600 116.060 ;
        RECT 32.535 113.700 33.055 115.690 ;
        RECT 31.990 112.090 33.600 113.700 ;
        RECT 32.535 110.100 33.055 112.090 ;
        RECT 31.990 108.490 33.600 110.100 ;
        RECT 32.535 106.500 33.055 108.490 ;
        RECT 25.115 105.545 29.335 106.185 ;
        RECT 20.820 105.310 21.180 105.340 ;
        RECT 20.130 105.010 21.180 105.310 ;
        RECT 25.115 105.275 26.220 105.545 ;
        RECT 20.820 104.980 21.180 105.010 ;
        RECT 31.990 104.890 33.600 106.500 ;
        RECT 32.535 102.900 33.055 104.890 ;
        RECT 31.990 101.290 33.600 102.900 ;
        RECT 32.535 99.300 33.055 101.290 ;
        RECT 31.990 97.690 33.600 99.300 ;
        RECT 32.535 95.700 33.055 97.690 ;
        RECT 31.990 94.090 33.600 95.700 ;
        RECT 32.535 92.100 33.055 94.090 ;
        RECT 31.990 90.490 33.600 92.100 ;
        RECT 32.535 88.500 33.055 90.490 ;
        RECT 31.990 86.890 33.600 88.500 ;
        RECT 32.535 85.895 33.055 86.890 ;
        RECT 34.935 85.895 35.455 118.295 ;
        RECT 9.125 73.700 27.960 74.220 ;
        RECT 27.535 70.140 27.960 73.700 ;
        RECT 27.400 69.580 28.085 70.140 ;
        RECT 27.550 63.225 28.240 63.780 ;
        RECT 27.650 62.205 28.175 63.225 ;
        RECT 27.650 61.445 28.180 62.205 ;
        RECT 38.590 61.445 39.110 120.420 ;
        RECT 44.585 89.515 44.885 217.610 ;
        RECT 46.565 122.425 46.865 218.900 ;
        RECT 46.315 121.625 47.120 122.425 ;
        RECT 44.310 88.715 45.115 89.515 ;
        RECT 49.000 70.220 50.500 220.760 ;
        RECT 62.870 213.670 63.170 224.760 ;
        RECT 66.575 220.820 66.875 224.760 ;
        RECT 70.215 224.760 70.230 224.890 ;
        RECT 84.935 224.760 84.950 224.900 ;
        RECT 88.605 224.760 88.630 225.130 ;
        RECT 92.610 224.760 92.615 225.030 ;
        RECT 96.290 224.760 96.295 224.875 ;
        RECT 107.010 224.760 107.030 224.940 ;
        RECT 110.700 224.760 110.710 224.850 ;
        RECT 114.385 224.760 114.390 224.940 ;
        RECT 118.370 224.760 118.375 225.210 ;
        RECT 70.215 220.860 70.515 224.760 ;
        RECT 84.935 222.940 85.235 224.760 ;
        RECT 88.605 222.955 88.905 224.760 ;
        RECT 84.840 222.455 85.360 222.940 ;
        RECT 88.500 222.470 89.020 222.955 ;
        RECT 66.560 220.490 66.890 220.820 ;
        RECT 70.200 220.530 70.530 220.860 ;
        RECT 62.775 213.235 63.355 213.670 ;
        RECT 92.315 210.930 92.615 224.760 ;
        RECT 52.825 210.630 92.615 210.930 ;
        RECT 48.990 68.440 50.510 70.220 ;
        RECT 27.650 60.925 39.110 61.445 ;
        RECT 28.685 59.465 29.310 59.605 ;
        RECT 4.210 59.155 29.310 59.465 ;
        RECT 28.685 59.095 29.310 59.155 ;
        RECT 28.690 59.090 29.305 59.095 ;
        RECT 22.730 57.270 23.980 57.440 ;
        RECT 13.360 56.370 23.980 57.270 ;
        RECT 0.995 35.135 1.000 36.290 ;
        RECT 2.500 35.135 2.505 36.290 ;
        RECT 2.500 23.170 2.510 25.490 ;
        RECT 13.360 7.720 14.260 56.370 ;
        RECT 22.730 56.360 23.980 56.370 ;
        RECT 23.060 48.560 25.760 50.500 ;
        RECT 13.370 5.770 14.260 7.720 ;
        RECT 23.930 7.480 24.830 48.560 ;
        RECT 23.925 6.740 24.830 7.480 ;
        RECT 33.990 3.560 34.890 59.725 ;
        RECT 49.000 5.000 50.500 68.440 ;
        RECT 52.825 64.910 53.125 210.630 ;
        RECT 95.995 209.710 96.295 224.760 ;
        RECT 54.150 209.410 96.295 209.710 ;
        RECT 54.150 65.650 54.450 209.410 ;
        RECT 99.670 208.775 99.970 224.760 ;
        RECT 54.960 208.475 99.970 208.775 ;
        RECT 54.960 66.400 55.260 208.475 ;
        RECT 103.350 207.980 103.650 224.760 ;
        RECT 55.820 207.680 103.650 207.980 ;
        RECT 55.820 67.220 56.120 207.680 ;
        RECT 107.010 206.980 107.310 224.760 ;
        RECT 56.640 206.680 107.310 206.980 ;
        RECT 56.640 67.950 56.940 206.680 ;
        RECT 110.700 206.135 111.000 224.760 ;
        RECT 57.620 205.835 111.000 206.135 ;
        RECT 57.620 68.860 57.920 205.835 ;
        RECT 114.385 205.205 114.685 224.760 ;
        RECT 58.710 204.905 114.685 205.205 ;
        RECT 58.710 69.565 59.010 204.905 ;
        RECT 118.075 204.225 118.375 224.760 ;
        RECT 59.735 203.925 118.375 204.225 ;
        RECT 121.740 224.760 121.750 224.960 ;
        RECT 128.945 224.760 129.110 225.415 ;
        RECT 129.410 224.760 129.545 225.415 ;
        RECT 59.735 70.340 60.035 203.925 ;
        RECT 121.740 203.040 122.040 224.760 ;
        RECT 61.010 202.740 122.040 203.040 ;
        RECT 61.010 71.205 61.310 202.740 ;
        RECT 125.430 197.760 125.730 224.760 ;
        RECT 67.335 197.460 125.730 197.760 ;
        RECT 67.335 189.360 67.635 197.460 ;
        RECT 67.320 189.030 67.650 189.360 ;
        RECT 76.485 147.950 78.085 194.670 ;
        RECT 79.785 147.950 81.385 194.670 ;
        RECT 88.560 147.950 90.160 194.670 ;
        RECT 91.860 147.950 93.460 194.670 ;
        RECT 100.635 147.950 102.235 194.670 ;
        RECT 103.935 147.950 105.535 194.670 ;
        RECT 112.710 147.950 114.310 194.670 ;
        RECT 116.010 147.950 117.610 194.670 ;
        RECT 128.945 189.635 129.545 224.760 ;
        RECT 132.540 224.760 132.790 225.360 ;
        RECT 133.090 224.760 133.140 225.360 ;
        RECT 128.940 189.025 129.550 189.635 ;
        RECT 132.540 154.275 133.140 224.760 ;
        RECT 136.320 224.760 136.470 225.400 ;
        RECT 136.770 224.760 136.920 225.400 ;
        RECT 136.320 215.770 136.920 224.760 ;
        RECT 139.980 224.760 140.150 225.360 ;
        RECT 140.450 224.760 140.580 225.360 ;
        RECT 139.980 217.440 140.580 224.760 ;
        RECT 143.660 224.760 143.830 225.340 ;
        RECT 144.130 224.760 144.260 225.340 ;
        RECT 143.660 219.620 144.260 224.760 ;
        RECT 147.350 224.760 147.510 225.265 ;
        RECT 147.810 224.760 147.950 225.265 ;
        RECT 151.490 224.760 152.660 225.585 ;
        RECT 147.350 221.455 147.950 224.760 ;
        RECT 147.320 220.845 147.980 221.455 ;
        RECT 143.605 218.905 144.325 219.620 ;
        RECT 139.920 216.725 140.640 217.440 ;
        RECT 136.265 215.055 136.985 215.770 ;
        RECT 132.535 153.665 133.145 154.275 ;
        RECT 80.935 140.035 81.835 140.075 ;
        RECT 80.195 138.950 81.835 140.035 ;
        RECT 78.590 124.050 80.430 125.685 ;
        RECT 61.010 70.905 71.645 71.205 ;
        RECT 59.735 70.040 70.185 70.340 ;
        RECT 58.710 69.265 68.980 69.565 ;
        RECT 57.620 68.560 68.025 68.860 ;
        RECT 56.640 67.650 67.070 67.950 ;
        RECT 55.820 66.920 66.045 67.220 ;
        RECT 54.960 66.100 65.060 66.400 ;
        RECT 54.150 65.350 64.060 65.650 ;
        RECT 52.825 64.610 62.840 64.910 ;
        RECT 53.130 8.675 54.030 61.775 ;
        RECT 53.125 7.780 54.035 8.675 ;
        RECT 33.990 2.660 46.910 3.560 ;
        RECT 46.010 1.000 46.910 2.660 ;
        RECT 53.130 1.870 54.030 7.780 ;
        RECT 55.390 3.875 56.290 57.505 ;
        RECT 62.540 9.500 62.840 64.610 ;
        RECT 63.760 10.270 64.060 65.350 ;
        RECT 64.760 11.335 65.060 66.100 ;
        RECT 65.745 12.100 66.045 66.920 ;
        RECT 66.770 12.885 67.070 67.650 ;
        RECT 67.725 13.480 68.025 68.560 ;
        RECT 68.680 14.150 68.980 69.265 ;
        RECT 69.885 15.045 70.185 70.040 ;
        RECT 71.345 16.015 71.645 70.905 ;
        RECT 71.150 15.215 71.955 16.015 ;
        RECT 69.770 14.560 70.290 15.045 ;
        RECT 68.575 13.665 69.095 14.150 ;
        RECT 67.610 12.995 68.130 13.480 ;
        RECT 66.655 12.400 67.175 12.885 ;
        RECT 65.625 11.615 66.145 12.100 ;
        RECT 64.650 10.850 65.170 11.335 ;
        RECT 63.640 9.785 64.160 10.270 ;
        RECT 62.440 9.015 62.960 9.500 ;
        RECT 79.050 4.550 79.950 124.050 ;
        RECT 80.935 6.480 81.835 138.950 ;
        RECT 82.960 139.050 111.080 139.950 ;
        RECT 82.960 8.415 83.860 139.050 ;
        RECT 152.060 135.880 152.660 224.760 ;
        RECT 154.870 224.045 155.170 224.760 ;
        RECT 154.280 222.745 156.080 224.045 ;
        RECT 155.965 218.935 156.615 219.590 ;
        RECT 153.605 217.380 154.255 217.405 ;
        RECT 153.605 216.780 155.510 217.380 ;
        RECT 153.605 216.750 154.255 216.780 ;
        RECT 153.840 215.090 154.490 215.745 ;
        RECT 152.030 135.270 152.690 135.880 ;
        RECT 153.865 89.585 154.465 215.090 ;
        RECT 97.905 28.860 99.505 89.180 ;
        RECT 101.205 28.860 102.805 89.180 ;
        RECT 113.200 28.860 114.800 89.180 ;
        RECT 116.500 28.860 118.100 89.180 ;
        RECT 128.495 28.860 130.095 89.180 ;
        RECT 131.795 28.860 133.395 89.180 ;
        RECT 143.790 28.860 145.390 89.180 ;
        RECT 147.090 28.860 148.690 89.180 ;
        RECT 153.860 88.975 154.470 89.585 ;
        RECT 154.910 69.185 155.510 216.780 ;
        RECT 154.905 68.575 155.515 69.185 ;
        RECT 155.980 48.785 156.580 218.935 ;
        RECT 155.975 48.175 156.585 48.785 ;
        RECT 157.225 28.415 157.825 221.425 ;
        RECT 157.200 27.750 157.855 28.415 ;
        RECT 82.960 7.515 157.310 8.415 ;
        RECT 80.935 5.580 135.230 6.480 ;
        RECT 55.390 2.975 75.970 3.875 ;
        RECT 79.050 3.650 113.150 4.550 ;
        RECT 75.070 2.430 75.970 2.975 ;
        RECT 53.130 1.000 68.990 1.870 ;
        RECT 75.070 1.530 91.070 2.430 ;
        RECT 90.170 1.000 91.070 1.530 ;
        RECT 112.250 1.000 113.150 3.650 ;
        RECT 134.330 1.000 135.230 5.580 ;
        RECT 156.410 1.000 157.310 7.515 ;
        RECT 53.130 0.970 68.090 1.000 ;
      LAYER via4 ;
        RECT 76.695 188.040 77.875 189.220 ;
        RECT 76.695 176.485 77.875 177.665 ;
        RECT 76.695 164.930 77.875 166.110 ;
        RECT 76.695 153.375 77.875 154.555 ;
        RECT 79.995 191.340 81.175 192.520 ;
        RECT 79.995 179.785 81.175 180.965 ;
        RECT 79.995 168.230 81.175 169.410 ;
        RECT 79.995 156.675 81.175 157.855 ;
        RECT 88.770 188.040 89.950 189.220 ;
        RECT 88.770 176.485 89.950 177.665 ;
        RECT 88.770 164.930 89.950 166.110 ;
        RECT 88.770 153.375 89.950 154.555 ;
        RECT 92.070 191.340 93.250 192.520 ;
        RECT 92.070 179.785 93.250 180.965 ;
        RECT 92.070 168.230 93.250 169.410 ;
        RECT 92.070 156.675 93.250 157.855 ;
        RECT 100.845 188.040 102.025 189.220 ;
        RECT 100.845 176.485 102.025 177.665 ;
        RECT 100.845 164.930 102.025 166.110 ;
        RECT 100.845 153.375 102.025 154.555 ;
        RECT 104.145 191.340 105.325 192.520 ;
        RECT 104.145 179.785 105.325 180.965 ;
        RECT 104.145 168.230 105.325 169.410 ;
        RECT 104.145 156.675 105.325 157.855 ;
        RECT 112.920 188.040 114.100 189.220 ;
        RECT 112.920 176.485 114.100 177.665 ;
        RECT 112.920 164.930 114.100 166.110 ;
        RECT 112.920 153.375 114.100 154.555 ;
        RECT 116.220 191.340 117.400 192.520 ;
        RECT 116.220 179.785 117.400 180.965 ;
        RECT 116.220 168.230 117.400 169.410 ;
        RECT 116.220 156.675 117.400 157.855 ;
        RECT 98.115 80.850 99.295 82.030 ;
        RECT 98.115 65.895 99.295 67.075 ;
        RECT 98.115 50.940 99.295 52.120 ;
        RECT 98.115 35.985 99.295 37.165 ;
        RECT 101.415 84.150 102.595 85.330 ;
        RECT 101.415 69.195 102.595 70.375 ;
        RECT 101.415 54.240 102.595 55.420 ;
        RECT 101.415 39.285 102.595 40.465 ;
        RECT 113.410 80.850 114.590 82.030 ;
        RECT 113.410 65.895 114.590 67.075 ;
        RECT 113.410 50.940 114.590 52.120 ;
        RECT 113.410 35.985 114.590 37.165 ;
        RECT 116.710 84.150 117.890 85.330 ;
        RECT 116.710 69.195 117.890 70.375 ;
        RECT 116.710 54.240 117.890 55.420 ;
        RECT 116.710 39.285 117.890 40.465 ;
        RECT 128.705 80.850 129.885 82.030 ;
        RECT 128.705 65.895 129.885 67.075 ;
        RECT 128.705 50.940 129.885 52.120 ;
        RECT 128.705 35.985 129.885 37.165 ;
        RECT 132.005 84.150 133.185 85.330 ;
        RECT 132.005 69.195 133.185 70.375 ;
        RECT 132.005 54.240 133.185 55.420 ;
        RECT 132.005 39.285 133.185 40.465 ;
        RECT 144.000 80.850 145.180 82.030 ;
        RECT 144.000 65.895 145.180 67.075 ;
        RECT 144.000 50.940 145.180 52.120 ;
        RECT 144.000 35.985 145.180 37.165 ;
        RECT 147.300 84.150 148.480 85.330 ;
        RECT 147.300 69.195 148.480 70.375 ;
        RECT 147.300 54.240 148.480 55.420 ;
        RECT 147.300 39.285 148.480 40.465 ;
      LAYER met5 ;
        RECT 71.010 191.130 119.790 192.730 ;
        RECT 71.010 187.830 119.790 189.430 ;
        RECT 71.010 179.575 119.790 181.175 ;
        RECT 71.010 176.275 119.790 177.875 ;
        RECT 71.010 168.020 119.790 169.620 ;
        RECT 71.010 164.720 119.790 166.320 ;
        RECT 71.010 156.465 119.790 158.065 ;
        RECT 71.010 153.165 119.790 154.765 ;
        RECT 90.820 83.940 152.480 85.540 ;
        RECT 90.820 80.640 152.480 82.240 ;
        RECT 90.820 68.985 152.480 70.585 ;
        RECT 90.820 65.685 152.480 67.285 ;
        RECT 90.820 54.030 152.480 55.630 ;
        RECT 90.820 50.730 152.480 52.330 ;
        RECT 90.820 39.075 152.480 40.675 ;
        RECT 90.820 35.775 152.480 37.375 ;
  END
END tt_um_mixed_signal_pulse_gen
END LIBRARY

