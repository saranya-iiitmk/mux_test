magic
tech sky130A
magscale 1 2
timestamp 1717180972
<< viali >>
rect 3249 11305 3283 11339
rect 9229 11305 9263 11339
rect 4629 11101 4663 11135
rect 3157 11033 3191 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 9137 11033 9171 11067
rect 4077 10965 4111 10999
rect 7297 10965 7331 10999
rect 2329 10761 2363 10795
rect 9045 10761 9079 10795
rect 5396 10693 5430 10727
rect 5733 10693 5767 10727
rect 1409 10625 1443 10659
rect 3065 10625 3099 10659
rect 3433 10625 3467 10659
rect 3617 10625 3651 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 10425 10625 10459 10659
rect 3341 10557 3375 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 7021 10557 7055 10591
rect 7113 10489 7147 10523
rect 1593 10421 1627 10455
rect 3525 10421 3559 10455
rect 4261 10421 4295 10455
rect 6377 10421 6411 10455
rect 10241 10421 10275 10455
rect 3341 10217 3375 10251
rect 3617 10217 3651 10251
rect 7665 10217 7699 10251
rect 8401 10217 8435 10251
rect 9413 10217 9447 10251
rect 8125 10149 8159 10183
rect 3341 10081 3375 10115
rect 3801 10081 3835 10115
rect 6285 10081 6319 10115
rect 8033 10081 8067 10115
rect 9597 10081 9631 10115
rect 2973 10013 3007 10047
rect 3430 10013 3464 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 9873 10013 9907 10047
rect 4046 9945 4080 9979
rect 5273 9945 5307 9979
rect 6552 9945 6586 9979
rect 7757 9945 7791 9979
rect 5181 9877 5215 9911
rect 6101 9877 6135 9911
rect 9689 9877 9723 9911
rect 6561 9673 6595 9707
rect 6745 9673 6779 9707
rect 7665 9673 7699 9707
rect 9312 9605 9346 9639
rect 3893 9537 3927 9571
rect 4169 9537 4203 9571
rect 6742 9537 6776 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 8309 9537 8343 9571
rect 8585 9537 8619 9571
rect 4813 9469 4847 9503
rect 5089 9469 5123 9503
rect 5641 9469 5675 9503
rect 7205 9469 7239 9503
rect 9045 9469 9079 9503
rect 7113 9401 7147 9435
rect 8401 9401 8435 9435
rect 3617 9333 3651 9367
rect 4077 9333 4111 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 8125 9333 8159 9367
rect 10425 9333 10459 9367
rect 4905 9129 4939 9163
rect 5641 9129 5675 9163
rect 4261 8993 4295 9027
rect 10425 8993 10459 9027
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 9689 8925 9723 8959
rect 9781 8925 9815 8959
rect 6377 8857 6411 8891
rect 7665 8857 7699 8891
rect 7849 8857 7883 8891
rect 8033 8857 8067 8891
rect 5825 8789 5859 8823
rect 9597 8789 9631 8823
rect 7113 8585 7147 8619
rect 6561 8517 6595 8551
rect 1593 8449 1627 8483
rect 4077 8449 4111 8483
rect 6745 8449 6779 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 7941 8449 7975 8483
rect 8208 8449 8242 8483
rect 1869 8381 1903 8415
rect 3341 8313 3375 8347
rect 3893 8245 3927 8279
rect 6377 8245 6411 8279
rect 9321 8245 9355 8279
rect 1593 8041 1627 8075
rect 6745 8041 6779 8075
rect 7113 8041 7147 8075
rect 9873 8041 9907 8075
rect 1869 7905 1903 7939
rect 3065 7905 3099 7939
rect 3525 7905 3559 7939
rect 9505 7905 9539 7939
rect 1961 7837 1995 7871
rect 3433 7837 3467 7871
rect 7665 7837 7699 7871
rect 8585 7837 8619 7871
rect 9321 7837 9355 7871
rect 9781 7837 9815 7871
rect 9965 7837 9999 7871
rect 10057 7837 10091 7871
rect 10241 7837 10275 7871
rect 5273 7769 5307 7803
rect 7941 7701 7975 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 10057 7701 10091 7735
rect 7757 7497 7791 7531
rect 8309 7497 8343 7531
rect 8677 7497 8711 7531
rect 9505 7497 9539 7531
rect 9413 7429 9447 7463
rect 10149 7429 10183 7463
rect 1685 7361 1719 7395
rect 3801 7361 3835 7395
rect 5917 7361 5951 7395
rect 6377 7361 6411 7395
rect 6633 7361 6667 7395
rect 8769 7361 8803 7395
rect 8953 7361 8987 7395
rect 10333 7361 10367 7395
rect 1961 7293 1995 7327
rect 4077 7293 4111 7327
rect 6193 7293 6227 7327
rect 8125 7293 8159 7327
rect 8217 7293 8251 7327
rect 9229 7293 9263 7327
rect 5733 7225 5767 7259
rect 3433 7157 3467 7191
rect 5549 7157 5583 7191
rect 6101 7157 6135 7191
rect 8953 7157 8987 7191
rect 9873 7157 9907 7191
rect 9965 7157 9999 7191
rect 1961 6953 1995 6987
rect 3985 6953 4019 6987
rect 8953 6953 8987 6987
rect 8769 6885 8803 6919
rect 2145 6817 2179 6851
rect 4997 6817 5031 6851
rect 5273 6817 5307 6851
rect 9505 6817 9539 6851
rect 10241 6817 10275 6851
rect 2237 6749 2271 6783
rect 3801 6749 3835 6783
rect 7389 6749 7423 6783
rect 5365 6681 5399 6715
rect 7634 6681 7668 6715
rect 6653 6613 6687 6647
rect 9689 6613 9723 6647
rect 7757 6409 7791 6443
rect 8953 6409 8987 6443
rect 10425 6409 10459 6443
rect 9290 6341 9324 6375
rect 3985 6273 4019 6307
rect 4629 6273 4663 6307
rect 6377 6273 6411 6307
rect 7941 6273 7975 6307
rect 8585 6273 8619 6307
rect 3893 6205 3927 6239
rect 4537 6205 4571 6239
rect 5089 6205 5123 6239
rect 8677 6205 8711 6239
rect 9045 6205 9079 6239
rect 4353 6137 4387 6171
rect 4997 6069 5031 6103
rect 5733 6069 5767 6103
rect 6561 6069 6595 6103
rect 1869 5865 1903 5899
rect 7297 5865 7331 5899
rect 8401 5865 8435 5899
rect 2421 5797 2455 5831
rect 2237 5729 2271 5763
rect 2881 5729 2915 5763
rect 3341 5729 3375 5763
rect 3617 5729 3651 5763
rect 4077 5729 4111 5763
rect 5825 5729 5859 5763
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 3249 5661 3283 5695
rect 5457 5661 5491 5695
rect 5549 5661 5583 5695
rect 8677 5661 8711 5695
rect 9781 5661 9815 5695
rect 9965 5661 9999 5695
rect 10149 5661 10183 5695
rect 4721 5525 4755 5559
rect 5273 5525 5307 5559
rect 8217 5525 8251 5559
rect 9229 5525 9263 5559
rect 9965 5525 9999 5559
rect 3985 5321 4019 5355
rect 5457 5253 5491 5287
rect 6653 5253 6687 5287
rect 8760 5253 8794 5287
rect 1961 5117 1995 5151
rect 2237 5117 2271 5151
rect 5733 5117 5767 5151
rect 6377 5117 6411 5151
rect 8493 5117 8527 5151
rect 3709 4981 3743 5015
rect 8125 4981 8159 5015
rect 9873 4981 9907 5015
rect 9229 4777 9263 4811
rect 9689 4777 9723 4811
rect 9321 4709 9355 4743
rect 4169 4641 4203 4675
rect 9137 4641 9171 4675
rect 10333 4641 10367 4675
rect 4445 4573 4479 4607
rect 7297 4573 7331 4607
rect 8033 4573 8067 4607
rect 8585 4573 8619 4607
rect 8953 4573 8987 4607
rect 9413 4573 9447 4607
rect 9781 4573 9815 4607
rect 7941 4437 7975 4471
rect 7205 4233 7239 4267
rect 8125 4233 8159 4267
rect 3341 4097 3375 4131
rect 4169 4097 4203 4131
rect 4629 4097 4663 4131
rect 7481 4097 7515 4131
rect 7573 4097 7607 4131
rect 7941 4097 7975 4131
rect 8769 4097 8803 4131
rect 9781 4097 9815 4131
rect 3433 4029 3467 4063
rect 3709 4029 3743 4063
rect 4077 4029 4111 4063
rect 4537 4029 4571 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 7665 4029 7699 4063
rect 8907 4029 8941 4063
rect 9045 4029 9079 4063
rect 9965 4029 9999 4063
rect 9321 3961 9355 3995
rect 3801 3893 3835 3927
rect 5825 3893 5859 3927
rect 7757 3893 7791 3927
rect 4537 3689 4571 3723
rect 5536 3689 5570 3723
rect 7021 3689 7055 3723
rect 8493 3689 8527 3723
rect 10425 3689 10459 3723
rect 8677 3621 8711 3655
rect 1593 3553 1627 3587
rect 5273 3553 5307 3587
rect 7113 3553 7147 3587
rect 9045 3553 9079 3587
rect 4353 3485 4387 3519
rect 5181 3485 5215 3519
rect 8769 3485 8803 3519
rect 1869 3417 1903 3451
rect 7380 3417 7414 3451
rect 9312 3417 9346 3451
rect 3341 3349 3375 3383
rect 3801 3349 3835 3383
rect 2421 3145 2455 3179
rect 9045 3145 9079 3179
rect 9873 3145 9907 3179
rect 10241 3145 10275 3179
rect 6193 3077 6227 3111
rect 7573 3077 7607 3111
rect 3525 3009 3559 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 7932 3009 7966 3043
rect 9229 3009 9263 3043
rect 10425 3009 10459 3043
rect 2973 2941 3007 2975
rect 3157 2941 3191 2975
rect 3617 2941 3651 2975
rect 7665 2941 7699 2975
rect 7297 2873 7331 2907
rect 4721 2805 4755 2839
rect 3065 2601 3099 2635
rect 5549 2601 5583 2635
rect 8033 2601 8067 2635
rect 9781 2601 9815 2635
rect 8401 2533 8435 2567
rect 3801 2465 3835 2499
rect 9505 2465 9539 2499
rect 10425 2465 10459 2499
rect 3249 2397 3283 2431
rect 7757 2397 7791 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 8493 2397 8527 2431
rect 8953 2397 8987 2431
rect 4077 2329 4111 2363
rect 7941 2261 7975 2295
<< metal1 >>
rect 1104 11450 10764 11472
rect 1104 11398 2157 11450
rect 2209 11398 2221 11450
rect 2273 11398 2285 11450
rect 2337 11398 2349 11450
rect 2401 11398 2413 11450
rect 2465 11398 4572 11450
rect 4624 11398 4636 11450
rect 4688 11398 4700 11450
rect 4752 11398 4764 11450
rect 4816 11398 4828 11450
rect 4880 11398 6987 11450
rect 7039 11398 7051 11450
rect 7103 11398 7115 11450
rect 7167 11398 7179 11450
rect 7231 11398 7243 11450
rect 7295 11398 9402 11450
rect 9454 11398 9466 11450
rect 9518 11398 9530 11450
rect 9582 11398 9594 11450
rect 9646 11398 9658 11450
rect 9710 11398 10764 11450
rect 1104 11376 10764 11398
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 3016 11308 3249 11336
rect 3016 11296 3022 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8996 11308 9229 11336
rect 8996 11296 9002 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3142 11024 3148 11076
rect 3200 11024 3206 11076
rect 6914 11024 6920 11076
rect 6972 11024 6978 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7374 11064 7380 11076
rect 7147 11036 7380 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 9122 11024 9128 11076
rect 9180 11024 9186 11076
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3384 10968 4077 10996
rect 3384 10956 3390 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4065 10959 4123 10965
rect 7285 10999 7343 11005
rect 7285 10965 7297 10999
rect 7331 10996 7343 10999
rect 8202 10996 8208 11008
rect 7331 10968 8208 10996
rect 7331 10965 7343 10968
rect 7285 10959 7343 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 1104 10906 10764 10928
rect 1104 10854 2817 10906
rect 2869 10854 2881 10906
rect 2933 10854 2945 10906
rect 2997 10854 3009 10906
rect 3061 10854 3073 10906
rect 3125 10854 5232 10906
rect 5284 10854 5296 10906
rect 5348 10854 5360 10906
rect 5412 10854 5424 10906
rect 5476 10854 5488 10906
rect 5540 10854 7647 10906
rect 7699 10854 7711 10906
rect 7763 10854 7775 10906
rect 7827 10854 7839 10906
rect 7891 10854 7903 10906
rect 7955 10854 10062 10906
rect 10114 10854 10126 10906
rect 10178 10854 10190 10906
rect 10242 10854 10254 10906
rect 10306 10854 10318 10906
rect 10370 10854 10764 10906
rect 1104 10832 10764 10854
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 3142 10792 3148 10804
rect 2363 10764 3148 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 8110 10792 8116 10804
rect 5920 10764 8116 10792
rect 5384 10727 5442 10733
rect 5384 10693 5396 10727
rect 5430 10724 5442 10727
rect 5721 10727 5779 10733
rect 5721 10724 5733 10727
rect 5430 10696 5733 10724
rect 5430 10693 5442 10696
rect 5384 10687 5442 10693
rect 5721 10693 5733 10696
rect 5767 10693 5779 10727
rect 5721 10687 5779 10693
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 5920 10665 5948 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9122 10792 9128 10804
rect 9079 10764 9128 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 8386 10724 8392 10736
rect 6012 10696 8392 10724
rect 6012 10665 6040 10696
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 5905 10659 5963 10665
rect 3651 10628 5764 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 4430 10588 4436 10600
rect 3375 10560 4436 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5736 10597 5764 10628
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6972 10628 7297 10656
rect 6972 10616 6978 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7742 10656 7748 10668
rect 7607 10628 7748 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8662 10656 8668 10668
rect 8343 10628 8668 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 3660 10492 4752 10520
rect 3660 10480 3666 10492
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3694 10452 3700 10464
rect 3559 10424 3700 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 4246 10412 4252 10464
rect 4304 10412 4310 10464
rect 4724 10452 4752 10492
rect 5644 10464 5672 10551
rect 5736 10520 5764 10551
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 5868 10560 7021 10588
rect 5868 10548 5874 10560
rect 7009 10557 7021 10560
rect 7055 10588 7067 10591
rect 7650 10588 7656 10600
rect 7055 10560 7656 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7101 10523 7159 10529
rect 7101 10520 7113 10523
rect 5736 10492 7113 10520
rect 7101 10489 7113 10492
rect 7147 10489 7159 10523
rect 7101 10483 7159 10489
rect 5626 10452 5632 10464
rect 4724 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 5776 10424 6377 10452
rect 5776 10412 5782 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8036 10452 8064 10619
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10459 10628 10916 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10888 10532 10916 10628
rect 10870 10480 10876 10532
rect 10928 10480 10934 10532
rect 7616 10424 8064 10452
rect 7616 10412 7622 10424
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9272 10424 10241 10452
rect 9272 10412 9278 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 1104 10362 10764 10384
rect 1104 10310 2157 10362
rect 2209 10310 2221 10362
rect 2273 10310 2285 10362
rect 2337 10310 2349 10362
rect 2401 10310 2413 10362
rect 2465 10310 4572 10362
rect 4624 10310 4636 10362
rect 4688 10310 4700 10362
rect 4752 10310 4764 10362
rect 4816 10310 4828 10362
rect 4880 10310 6987 10362
rect 7039 10310 7051 10362
rect 7103 10310 7115 10362
rect 7167 10310 7179 10362
rect 7231 10310 7243 10362
rect 7295 10310 9402 10362
rect 9454 10310 9466 10362
rect 9518 10310 9530 10362
rect 9582 10310 9594 10362
rect 9646 10310 9658 10362
rect 9710 10310 10764 10362
rect 1104 10288 10764 10310
rect 1578 10208 1584 10260
rect 1636 10208 1642 10260
rect 3326 10208 3332 10260
rect 3384 10208 3390 10260
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3476 10220 3617 10248
rect 3476 10208 3482 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 5718 10248 5724 10260
rect 3605 10211 3663 10217
rect 3804 10220 5724 10248
rect 1596 10044 1624 10208
rect 3804 10180 3832 10220
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 8386 10208 8392 10260
rect 8444 10208 8450 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 10686 10248 10692 10260
rect 9447 10220 10692 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 3344 10152 3832 10180
rect 3344 10121 3372 10152
rect 8110 10140 8116 10192
rect 8168 10140 8174 10192
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 1596 10016 2973 10044
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3418 10047 3476 10053
rect 3418 10013 3430 10047
rect 3464 10046 3476 10047
rect 3464 10018 3556 10046
rect 3464 10013 3476 10018
rect 3418 10007 3476 10013
rect 3528 9908 3556 10018
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3804 10044 3832 10075
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5684 10084 6285 10112
rect 5684 10072 5690 10084
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 7742 10072 7748 10124
rect 7800 10072 7806 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8478 10112 8484 10124
rect 8067 10084 8484 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 3660 10016 3832 10044
rect 3660 10004 3666 10016
rect 5810 10004 5816 10056
rect 5868 10004 5874 10056
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10044 6055 10047
rect 6822 10044 6828 10056
rect 6043 10016 6828 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 3694 9936 3700 9988
rect 3752 9976 3758 9988
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 3752 9948 4046 9976
rect 3752 9936 3758 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 4034 9939 4092 9945
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 4764 9948 5273 9976
rect 4764 9936 4770 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 5261 9939 5319 9945
rect 3878 9908 3884 9920
rect 3528 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9908 3942 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 3936 9880 5181 9908
rect 3936 9868 3942 9880
rect 5169 9877 5181 9880
rect 5215 9908 5227 9911
rect 6012 9908 6040 10007
rect 6822 10004 6828 10016
rect 6880 10044 6886 10056
rect 7760 10044 7788 10072
rect 6880 10016 7788 10044
rect 7929 10047 7987 10053
rect 6880 10004 6886 10016
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 6546 9985 6552 9988
rect 6540 9939 6552 9985
rect 6546 9936 6552 9939
rect 6604 9936 6610 9988
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7745 9979 7803 9985
rect 7745 9976 7757 9979
rect 7156 9948 7757 9976
rect 7156 9936 7162 9948
rect 7745 9945 7757 9948
rect 7791 9945 7803 9979
rect 7944 9976 7972 10007
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 8404 10053 8432 10084
rect 8478 10072 8484 10084
rect 8536 10112 8542 10124
rect 9214 10112 9220 10124
rect 8536 10084 9220 10112
rect 8536 10072 8542 10084
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9232 10044 9260 10072
rect 9171 10016 9260 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 8588 9976 8616 10007
rect 9416 9976 9444 10211
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9631 10084 9904 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9876 10053 9904 10084
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 7944 9948 9444 9976
rect 7745 9939 7803 9945
rect 5215 9880 6040 9908
rect 6089 9911 6147 9917
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 7374 9908 7380 9920
rect 6135 9880 7380 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9548 9880 9689 9908
rect 9548 9868 9554 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 1104 9818 10764 9840
rect 1104 9766 2817 9818
rect 2869 9766 2881 9818
rect 2933 9766 2945 9818
rect 2997 9766 3009 9818
rect 3061 9766 3073 9818
rect 3125 9766 5232 9818
rect 5284 9766 5296 9818
rect 5348 9766 5360 9818
rect 5412 9766 5424 9818
rect 5476 9766 5488 9818
rect 5540 9766 7647 9818
rect 7699 9766 7711 9818
rect 7763 9766 7775 9818
rect 7827 9766 7839 9818
rect 7891 9766 7903 9818
rect 7955 9766 10062 9818
rect 10114 9766 10126 9818
rect 10178 9766 10190 9818
rect 10242 9766 10254 9818
rect 10306 9766 10318 9818
rect 10370 9766 10764 9818
rect 1104 9744 10764 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3602 9704 3608 9716
rect 2740 9676 3608 9704
rect 2740 9664 2746 9676
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 4706 9664 4712 9716
rect 4764 9664 4770 9716
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6696 9676 6745 9704
rect 6696 9664 6702 9676
rect 6733 9673 6745 9676
rect 6779 9704 6791 9707
rect 7558 9704 7564 9716
rect 6779 9676 7564 9704
rect 6779 9673 6791 9676
rect 6733 9667 6791 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7653 9707 7711 9713
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 8110 9704 8116 9716
rect 7699 9676 8116 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8478 9664 8484 9716
rect 8536 9664 8542 9716
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4724 9568 4752 9664
rect 5736 9608 7328 9636
rect 5736 9580 5764 9608
rect 4203 9540 4752 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 6730 9571 6788 9577
rect 6730 9537 6742 9571
rect 6776 9568 6788 9571
rect 7098 9568 7104 9580
rect 6776 9540 7104 9568
rect 6776 9537 6788 9540
rect 6730 9531 6788 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7300 9577 7328 9608
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8496 9568 8524 9664
rect 9300 9639 9358 9645
rect 9300 9605 9312 9639
rect 9346 9636 9358 9639
rect 9490 9636 9496 9648
rect 9346 9608 9496 9636
rect 9346 9605 9358 9608
rect 9300 9599 9358 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8343 9540 8432 9568
rect 8496 9540 8585 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4488 9472 4813 9500
rect 4488 9460 4494 9472
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 6914 9500 6920 9512
rect 5675 9472 6920 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7484 9500 7512 9528
rect 7239 9472 7512 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 8110 9460 8116 9512
rect 8168 9460 8174 9512
rect 4246 9432 4252 9444
rect 4080 9404 4252 9432
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 4080 9373 4108 9404
rect 4246 9392 4252 9404
rect 4304 9432 4310 9444
rect 5442 9432 5448 9444
rect 4304 9404 5448 9432
rect 4304 9392 4310 9404
rect 5442 9392 5448 9404
rect 5500 9432 5506 9444
rect 7101 9435 7159 9441
rect 5500 9404 6316 9432
rect 5500 9392 5506 9404
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6052 9336 6193 9364
rect 6052 9324 6058 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6288 9364 6316 9404
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 8128 9432 8156 9460
rect 8404 9441 8432 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9030 9460 9036 9512
rect 9088 9460 9094 9512
rect 7147 9404 8156 9432
rect 8389 9435 8447 9441
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 8389 9401 8401 9435
rect 8435 9401 8447 9435
rect 8389 9395 8447 9401
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6288 9336 7297 9364
rect 6181 9327 6239 9333
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8202 9364 8208 9376
rect 8159 9336 8208 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10459 9336 10824 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 1104 9274 10764 9296
rect 1104 9222 2157 9274
rect 2209 9222 2221 9274
rect 2273 9222 2285 9274
rect 2337 9222 2349 9274
rect 2401 9222 2413 9274
rect 2465 9222 4572 9274
rect 4624 9222 4636 9274
rect 4688 9222 4700 9274
rect 4752 9222 4764 9274
rect 4816 9222 4828 9274
rect 4880 9222 6987 9274
rect 7039 9222 7051 9274
rect 7103 9222 7115 9274
rect 7167 9222 7179 9274
rect 7231 9222 7243 9274
rect 7295 9222 9402 9274
rect 9454 9222 9466 9274
rect 9518 9222 9530 9274
rect 9582 9222 9594 9274
rect 9646 9222 9658 9274
rect 9710 9222 10764 9274
rect 1104 9200 10764 9222
rect 3602 9120 3608 9172
rect 3660 9120 3666 9172
rect 4430 9120 4436 9172
rect 4488 9120 4494 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5074 9160 5080 9172
rect 4939 9132 5080 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 5718 9160 5724 9172
rect 5675 9132 5724 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 3620 9024 3648 9120
rect 4448 9092 4476 9120
rect 6638 9092 6644 9104
rect 4448 9064 6644 9092
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 3620 8996 4261 9024
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 5442 8956 5448 8968
rect 5399 8928 5448 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6196 8965 6224 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10796 9024 10824 9336
rect 10459 8996 10824 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9723 8928 9781 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6365 8891 6423 8897
rect 6365 8888 6377 8891
rect 5684 8860 6377 8888
rect 5684 8848 5690 8860
rect 6365 8857 6377 8860
rect 6411 8857 6423 8891
rect 6365 8851 6423 8857
rect 7374 8848 7380 8900
rect 7432 8888 7438 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7432 8860 7665 8888
rect 7432 8848 7438 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 7837 8891 7895 8897
rect 7837 8857 7849 8891
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 6914 8820 6920 8832
rect 5859 8792 6920 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7852 8820 7880 8851
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 9858 8888 9864 8900
rect 8076 8860 9864 8888
rect 8076 8848 8082 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 8110 8820 8116 8832
rect 7852 8792 8116 8820
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 9214 8780 9220 8832
rect 9272 8820 9278 8832
rect 9585 8823 9643 8829
rect 9585 8820 9597 8823
rect 9272 8792 9597 8820
rect 9272 8780 9278 8792
rect 9585 8789 9597 8792
rect 9631 8789 9643 8823
rect 9585 8783 9643 8789
rect 1104 8730 10764 8752
rect 1104 8678 2817 8730
rect 2869 8678 2881 8730
rect 2933 8678 2945 8730
rect 2997 8678 3009 8730
rect 3061 8678 3073 8730
rect 3125 8678 5232 8730
rect 5284 8678 5296 8730
rect 5348 8678 5360 8730
rect 5412 8678 5424 8730
rect 5476 8678 5488 8730
rect 5540 8678 7647 8730
rect 7699 8678 7711 8730
rect 7763 8678 7775 8730
rect 7827 8678 7839 8730
rect 7891 8678 7903 8730
rect 7955 8678 10062 8730
rect 10114 8678 10126 8730
rect 10178 8678 10190 8730
rect 10242 8678 10254 8730
rect 10306 8678 10318 8730
rect 10370 8678 10764 8730
rect 1104 8656 10764 8678
rect 6730 8616 6736 8628
rect 6564 8588 6736 8616
rect 6564 8557 6592 8588
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 8386 8616 8392 8628
rect 7147 8588 8392 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 6549 8551 6607 8557
rect 6549 8517 6561 8551
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 3326 8480 3332 8492
rect 2990 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3988 8452 4077 8480
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 3988 8356 4016 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 6564 8412 6592 8511
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 9048 8548 9076 8576
rect 6880 8520 9076 8548
rect 6880 8508 6886 8520
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6914 8480 6920 8492
rect 6779 8452 6920 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 7944 8489 7972 8520
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6972 8452 7297 8480
rect 6972 8440 6978 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 7484 8412 7512 8443
rect 6564 8384 7512 8412
rect 7576 8412 7604 8443
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8202 8489 8208 8492
rect 8196 8480 8208 8489
rect 8163 8452 8208 8480
rect 8196 8443 8208 8452
rect 8202 8440 8208 8443
rect 8260 8440 8266 8492
rect 8036 8412 8064 8440
rect 7576 8384 8064 8412
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 3970 8344 3976 8356
rect 3375 8316 3976 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 3878 8236 3884 8288
rect 3936 8236 3942 8288
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6328 8248 6377 8276
rect 6328 8236 6334 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6365 8239 6423 8245
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 1104 8186 10764 8208
rect 1104 8134 2157 8186
rect 2209 8134 2221 8186
rect 2273 8134 2285 8186
rect 2337 8134 2349 8186
rect 2401 8134 2413 8186
rect 2465 8134 4572 8186
rect 4624 8134 4636 8186
rect 4688 8134 4700 8186
rect 4752 8134 4764 8186
rect 4816 8134 4828 8186
rect 4880 8134 6987 8186
rect 7039 8134 7051 8186
rect 7103 8134 7115 8186
rect 7167 8134 7179 8186
rect 7231 8134 7243 8186
rect 7295 8134 9402 8186
rect 9454 8134 9466 8186
rect 9518 8134 9530 8186
rect 9582 8134 9594 8186
rect 9646 8134 9658 8186
rect 9710 8134 10764 8186
rect 1104 8112 10764 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1854 8072 1860 8084
rect 1627 8044 1860 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 6822 8072 6828 8084
rect 6779 8044 6828 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7466 8072 7472 8084
rect 7147 8044 7472 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 6086 7964 6092 8016
rect 6144 8004 6150 8016
rect 7116 8004 7144 8035
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 9858 8032 9864 8084
rect 9916 8032 9922 8084
rect 6144 7976 7144 8004
rect 6144 7964 6150 7976
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7905 1915 7939
rect 1857 7899 1915 7905
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3142 7936 3148 7948
rect 3099 7908 3148 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 1872 7800 1900 7899
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3344 7908 3525 7936
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 3344 7868 3372 7908
rect 3513 7905 3525 7908
rect 3559 7936 3571 7939
rect 3878 7936 3884 7948
rect 3559 7908 3884 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 9122 7936 9128 7948
rect 6288 7908 9128 7936
rect 6288 7880 6316 7908
rect 9122 7896 9128 7908
rect 9180 7936 9186 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9180 7908 9505 7936
rect 9180 7896 9186 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 10594 7936 10600 7948
rect 9493 7899 9551 7905
rect 9968 7908 10600 7936
rect 1995 7840 3372 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7616 7840 7665 7868
rect 7616 7828 7622 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9968 7877 9996 7908
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 9953 7871 10011 7877
rect 9815 7840 9904 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 3602 7800 3608 7812
rect 1872 7772 3608 7800
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 6178 7800 6184 7812
rect 5307 7772 6184 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 9876 7744 9904 7840
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10275 7840 10824 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10060 7800 10088 7831
rect 10060 7772 10456 7800
rect 10428 7744 10456 7772
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8018 7732 8024 7744
rect 7975 7704 8024 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8352 7704 8953 7732
rect 8352 7692 8358 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9766 7732 9772 7744
rect 9447 7704 9772 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 9858 7692 9864 7744
rect 9916 7692 9922 7744
rect 9950 7692 9956 7744
rect 10008 7732 10014 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 10008 7704 10057 7732
rect 10008 7692 10014 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 1104 7642 10764 7664
rect 1104 7590 2817 7642
rect 2869 7590 2881 7642
rect 2933 7590 2945 7642
rect 2997 7590 3009 7642
rect 3061 7590 3073 7642
rect 3125 7590 5232 7642
rect 5284 7590 5296 7642
rect 5348 7590 5360 7642
rect 5412 7590 5424 7642
rect 5476 7590 5488 7642
rect 5540 7590 7647 7642
rect 7699 7590 7711 7642
rect 7763 7590 7775 7642
rect 7827 7590 7839 7642
rect 7891 7590 7903 7642
rect 7955 7590 10062 7642
rect 10114 7590 10126 7642
rect 10178 7590 10190 7642
rect 10242 7590 10254 7642
rect 10306 7590 10318 7642
rect 10370 7590 10764 7642
rect 1104 7568 10764 7590
rect 2682 7528 2688 7540
rect 1688 7500 2688 7528
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1688 7401 1716 7500
rect 2682 7488 2688 7500
rect 2740 7528 2746 7540
rect 2740 7500 6408 7528
rect 2740 7488 2746 7500
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 3326 7392 3332 7404
rect 3082 7378 3332 7392
rect 1673 7355 1731 7361
rect 3068 7364 3332 7378
rect 1946 7284 1952 7336
rect 2004 7284 2010 7336
rect 3068 7256 3096 7364
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3804 7401 3832 7500
rect 6380 7460 6408 7500
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7616 7500 7757 7528
rect 7616 7488 7622 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 8294 7488 8300 7540
rect 8352 7488 8358 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 8665 7531 8723 7537
rect 8665 7528 8677 7531
rect 8628 7500 8677 7528
rect 8628 7488 8634 7500
rect 8665 7497 8677 7500
rect 8711 7497 8723 7531
rect 8665 7491 8723 7497
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 9272 7500 9505 7528
rect 9272 7488 9278 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 9493 7491 9551 7497
rect 6840 7460 6868 7488
rect 6380 7432 6868 7460
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 5626 7392 5632 7404
rect 5198 7378 5632 7392
rect 3789 7355 3847 7361
rect 5184 7364 5632 7378
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3200 7296 4077 7324
rect 3200 7284 3206 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 3068 7228 3556 7256
rect 3418 7148 3424 7200
rect 3476 7148 3482 7200
rect 3528 7188 3556 7228
rect 5184 7188 5212 7364
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6270 7392 6276 7404
rect 5951 7364 6276 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6380 7401 6408 7432
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9401 7463 9459 7469
rect 8168 7432 8800 7460
rect 8168 7420 8174 7432
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 6365 7355 6423 7361
rect 6472 7364 6633 7392
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 6144 7296 6193 7324
rect 6144 7284 6150 7296
rect 6181 7293 6193 7296
rect 6227 7293 6239 7327
rect 6472 7324 6500 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 8386 7392 8392 7404
rect 6621 7355 6679 7361
rect 8128 7364 8392 7392
rect 8128 7333 8156 7364
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8772 7401 8800 7432
rect 9401 7429 9413 7463
rect 9447 7460 9459 7463
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9447 7432 10149 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 10137 7429 10149 7432
rect 10183 7460 10195 7463
rect 10183 7432 10456 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10428 7404 10456 7432
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 8987 7364 9904 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9876 7336 9904 7364
rect 10318 7352 10324 7404
rect 10376 7352 10382 7404
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 6181 7287 6239 7293
rect 6380 7296 6500 7324
rect 8113 7327 8171 7333
rect 5721 7259 5779 7265
rect 5721 7225 5733 7259
rect 5767 7256 5779 7259
rect 6380 7256 6408 7296
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 8570 7324 8576 7336
rect 8251 7296 8576 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9180 7296 9229 7324
rect 9180 7284 9186 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10336 7324 10364 7352
rect 10796 7324 10824 7840
rect 9916 7296 9996 7324
rect 10336 7296 10824 7324
rect 9916 7284 9922 7296
rect 5767 7228 6408 7256
rect 5767 7225 5779 7228
rect 5721 7219 5779 7225
rect 3528 7160 5212 7188
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 6135 7160 8953 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 8941 7157 8953 7160
rect 8987 7157 8999 7191
rect 8941 7151 8999 7157
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 9968 7197 9996 7296
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7188 10011 7191
rect 10502 7188 10508 7200
rect 9999 7160 10508 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 1104 7098 10764 7120
rect 1104 7046 2157 7098
rect 2209 7046 2221 7098
rect 2273 7046 2285 7098
rect 2337 7046 2349 7098
rect 2401 7046 2413 7098
rect 2465 7046 4572 7098
rect 4624 7046 4636 7098
rect 4688 7046 4700 7098
rect 4752 7046 4764 7098
rect 4816 7046 4828 7098
rect 4880 7046 6987 7098
rect 7039 7046 7051 7098
rect 7103 7046 7115 7098
rect 7167 7046 7179 7098
rect 7231 7046 7243 7098
rect 7295 7046 9402 7098
rect 9454 7046 9466 7098
rect 9518 7046 9530 7098
rect 9582 7046 9594 7098
rect 9646 7046 9658 7098
rect 9710 7046 10764 7098
rect 1104 7024 10764 7046
rect 1946 6944 1952 6996
rect 2004 6944 2010 6996
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 3660 6956 3985 6984
rect 3660 6944 3666 6956
rect 3973 6953 3985 6956
rect 4019 6953 4031 6987
rect 3973 6947 4031 6953
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 10318 6916 10324 6928
rect 8803 6888 10324 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 1912 6820 2145 6848
rect 1912 6808 1918 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 3142 6848 3148 6860
rect 2133 6811 2191 6817
rect 2746 6820 3148 6848
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2746 6780 2774 6820
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 3384 6820 4997 6848
rect 3384 6808 3390 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5534 6848 5540 6860
rect 5307 6820 5540 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 9508 6857 9536 6888
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 9916 6820 10241 6848
rect 9916 6808 9922 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 3418 6780 3424 6792
rect 2271 6752 2774 6780
rect 3160 6752 3424 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 3160 6656 3188 6752
rect 3418 6740 3424 6752
rect 3476 6780 3482 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3476 6752 3801 6780
rect 3476 6740 3482 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7423 6752 8524 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4212 6684 5365 6712
rect 4212 6672 4218 6684
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 7622 6715 7680 6721
rect 7622 6712 7634 6715
rect 7524 6684 7634 6712
rect 7524 6672 7530 6684
rect 7622 6681 7634 6684
rect 7668 6681 7680 6715
rect 7622 6675 7680 6681
rect 8496 6656 8524 6752
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6236 6616 6653 6644
rect 6236 6604 6242 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 8478 6604 8484 6656
rect 8536 6604 8542 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 1104 6554 10764 6576
rect 1104 6502 2817 6554
rect 2869 6502 2881 6554
rect 2933 6502 2945 6554
rect 2997 6502 3009 6554
rect 3061 6502 3073 6554
rect 3125 6502 5232 6554
rect 5284 6502 5296 6554
rect 5348 6502 5360 6554
rect 5412 6502 5424 6554
rect 5476 6502 5488 6554
rect 5540 6502 7647 6554
rect 7699 6502 7711 6554
rect 7763 6502 7775 6554
rect 7827 6502 7839 6554
rect 7891 6502 7903 6554
rect 7955 6502 10062 6554
rect 10114 6502 10126 6554
rect 10178 6502 10190 6554
rect 10242 6502 10254 6554
rect 10306 6502 10318 6554
rect 10370 6502 10764 6554
rect 1104 6480 10764 6502
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7745 6443 7803 6449
rect 7745 6440 7757 6443
rect 7524 6412 7757 6440
rect 7524 6400 7530 6412
rect 7745 6409 7757 6412
rect 7791 6409 7803 6443
rect 7745 6403 7803 6409
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 4890 6304 4896 6316
rect 4663 6276 4896 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5684 6276 6377 6304
rect 5684 6264 5690 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8036 6304 8064 6400
rect 8956 6372 8984 6403
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 9278 6375 9336 6381
rect 9278 6372 9290 6375
rect 8956 6344 9290 6372
rect 9278 6341 9290 6344
rect 9324 6341 9336 6375
rect 9278 6335 9336 6341
rect 7975 6276 8064 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8444 6276 8585 6304
rect 8444 6264 8450 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 9692 6304 9720 6400
rect 8573 6267 8631 6273
rect 8680 6276 9720 6304
rect 3326 6196 3332 6248
rect 3384 6196 3390 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 8680 6245 8708 6276
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3660 6208 3893 6236
rect 3660 6196 3666 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 3881 6199 3939 6205
rect 4172 6208 4537 6236
rect 3344 6168 3372 6196
rect 4172 6168 4200 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 3344 6140 4200 6168
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 5092 6168 5120 6199
rect 9048 6168 9076 6199
rect 4387 6140 5120 6168
rect 8496 6140 9076 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 8496 6112 8524 6140
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5626 6100 5632 6112
rect 5031 6072 5632 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 6052 6072 6561 6100
rect 6052 6060 6058 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 1104 6010 10764 6032
rect 1104 5958 2157 6010
rect 2209 5958 2221 6010
rect 2273 5958 2285 6010
rect 2337 5958 2349 6010
rect 2401 5958 2413 6010
rect 2465 5958 4572 6010
rect 4624 5958 4636 6010
rect 4688 5958 4700 6010
rect 4752 5958 4764 6010
rect 4816 5958 4828 6010
rect 4880 5958 6987 6010
rect 7039 5958 7051 6010
rect 7103 5958 7115 6010
rect 7167 5958 7179 6010
rect 7231 5958 7243 6010
rect 7295 5958 9402 6010
rect 9454 5958 9466 6010
rect 9518 5958 9530 6010
rect 9582 5958 9594 6010
rect 9646 5958 9658 6010
rect 9710 5958 10764 6010
rect 1104 5936 10764 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 8110 5896 8116 5908
rect 7331 5868 8116 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 8110 5856 8116 5868
rect 8168 5896 8174 5908
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 8168 5868 8401 5896
rect 8168 5856 8174 5868
rect 8389 5865 8401 5868
rect 8435 5865 8447 5899
rect 8389 5859 8447 5865
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5797 2467 5831
rect 2409 5791 2467 5797
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2424 5760 2452 5791
rect 2271 5732 2452 5760
rect 2869 5763 2927 5769
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 3142 5760 3148 5772
rect 2915 5732 3148 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 3326 5720 3332 5772
rect 3384 5720 3390 5772
rect 3605 5763 3663 5769
rect 3605 5729 3617 5763
rect 3651 5760 3663 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3651 5732 4077 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 9968 5760 9996 5856
rect 9968 5732 10180 5760
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2777 5695 2835 5701
rect 2179 5664 2268 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2240 5568 2268 5664
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3050 5692 3056 5704
rect 2823 5664 3056 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3970 5692 3976 5704
rect 3283 5664 3976 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3970 5652 3976 5664
rect 4028 5692 4034 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4028 5664 5457 5692
rect 4028 5652 4034 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 8711 5664 8984 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 5552 5624 5580 5655
rect 5552 5596 5672 5624
rect 5644 5568 5672 5596
rect 6012 5596 6302 5624
rect 6012 5568 6040 5596
rect 8956 5568 8984 5664
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 10152 5701 10180 5732
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 9968 5624 9996 5655
rect 10502 5624 10508 5636
rect 9968 5596 10508 5624
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 2222 5516 2228 5568
rect 2280 5516 2286 5568
rect 4706 5516 4712 5568
rect 4764 5516 4770 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4948 5528 5273 5556
rect 4948 5516 4954 5528
rect 5261 5525 5273 5528
rect 5307 5525 5319 5559
rect 5261 5519 5319 5525
rect 5626 5516 5632 5568
rect 5684 5516 5690 5568
rect 5994 5516 6000 5568
rect 6052 5516 6058 5568
rect 8202 5516 8208 5568
rect 8260 5516 8266 5568
rect 8938 5516 8944 5568
rect 8996 5516 9002 5568
rect 9214 5516 9220 5568
rect 9272 5516 9278 5568
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 9916 5528 9965 5556
rect 9916 5516 9922 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 1104 5466 10764 5488
rect 1104 5414 2817 5466
rect 2869 5414 2881 5466
rect 2933 5414 2945 5466
rect 2997 5414 3009 5466
rect 3061 5414 3073 5466
rect 3125 5414 5232 5466
rect 5284 5414 5296 5466
rect 5348 5414 5360 5466
rect 5412 5414 5424 5466
rect 5476 5414 5488 5466
rect 5540 5414 7647 5466
rect 7699 5414 7711 5466
rect 7763 5414 7775 5466
rect 7827 5414 7839 5466
rect 7891 5414 7903 5466
rect 7955 5414 10062 5466
rect 10114 5414 10126 5466
rect 10178 5414 10190 5466
rect 10242 5414 10254 5466
rect 10306 5414 10318 5466
rect 10370 5414 10764 5466
rect 1104 5392 10764 5414
rect 3970 5312 3976 5364
rect 4028 5312 4034 5364
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 4764 5324 5488 5352
rect 4764 5312 4770 5324
rect 5460 5293 5488 5324
rect 5994 5312 6000 5364
rect 6052 5352 6058 5364
rect 6052 5324 6776 5352
rect 6052 5312 6058 5324
rect 5445 5287 5503 5293
rect 5445 5253 5457 5287
rect 5491 5253 5503 5287
rect 5445 5247 5503 5253
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 5776 5256 6653 5284
rect 5776 5244 5782 5256
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 6748 5284 6776 5324
rect 8748 5287 8806 5293
rect 6748 5256 7130 5284
rect 6641 5247 6699 5253
rect 8748 5253 8760 5287
rect 8794 5284 8806 5287
rect 9214 5284 9220 5296
rect 8794 5256 9220 5284
rect 8794 5253 8806 5256
rect 8748 5247 8806 5253
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 3358 5188 4370 5216
rect 1946 5108 1952 5160
rect 2004 5108 2010 5160
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 2682 5148 2688 5160
rect 2280 5120 2688 5148
rect 2280 5108 2286 5120
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3436 5024 3464 5188
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5644 5120 5733 5148
rect 5644 5024 5672 5120
rect 5721 5117 5733 5120
rect 5767 5148 5779 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5767 5120 6377 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 8478 5108 8484 5160
rect 8536 5108 8542 5160
rect 3418 4972 3424 5024
rect 3476 4972 3482 5024
rect 3694 4972 3700 5024
rect 3752 4972 3758 5024
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8754 5012 8760 5024
rect 8159 4984 8760 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9858 4972 9864 5024
rect 9916 4972 9922 5024
rect 1104 4922 10764 4944
rect 1104 4870 2157 4922
rect 2209 4870 2221 4922
rect 2273 4870 2285 4922
rect 2337 4870 2349 4922
rect 2401 4870 2413 4922
rect 2465 4870 4572 4922
rect 4624 4870 4636 4922
rect 4688 4870 4700 4922
rect 4752 4870 4764 4922
rect 4816 4870 4828 4922
rect 4880 4870 6987 4922
rect 7039 4870 7051 4922
rect 7103 4870 7115 4922
rect 7167 4870 7179 4922
rect 7231 4870 7243 4922
rect 7295 4870 9402 4922
rect 9454 4870 9466 4922
rect 9518 4870 9530 4922
rect 9582 4870 9594 4922
rect 9646 4870 9658 4922
rect 9710 4870 10764 4922
rect 1104 4848 10764 4870
rect 3694 4768 3700 4820
rect 3752 4768 3758 4820
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 8168 4780 9229 4808
rect 8168 4768 8174 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9766 4808 9772 4820
rect 9723 4780 9772 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 3712 4672 3740 4768
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 9309 4743 9367 4749
rect 9309 4740 9321 4743
rect 7432 4712 9321 4740
rect 7432 4700 7438 4712
rect 9309 4709 9321 4712
rect 9355 4709 9367 4743
rect 9309 4703 9367 4709
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 3712 4644 4169 4672
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 4157 4635 4215 4641
rect 8772 4644 9137 4672
rect 8772 4616 8800 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9916 4644 10333 4672
rect 9916 4632 9922 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4448 4480 4476 4567
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7524 4576 8033 4604
rect 7524 4564 7530 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8570 4564 8576 4616
rect 8628 4564 8634 4616
rect 8754 4564 8760 4616
rect 8812 4564 8818 4616
rect 8938 4564 8944 4616
rect 8996 4564 9002 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9447 4576 9781 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7616 4440 7941 4468
rect 7616 4428 7622 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 1104 4378 10764 4400
rect 1104 4326 2817 4378
rect 2869 4326 2881 4378
rect 2933 4326 2945 4378
rect 2997 4326 3009 4378
rect 3061 4326 3073 4378
rect 3125 4326 5232 4378
rect 5284 4326 5296 4378
rect 5348 4326 5360 4378
rect 5412 4326 5424 4378
rect 5476 4326 5488 4378
rect 5540 4326 7647 4378
rect 7699 4326 7711 4378
rect 7763 4326 7775 4378
rect 7827 4326 7839 4378
rect 7891 4326 7903 4378
rect 7955 4326 10062 4378
rect 10114 4326 10126 4378
rect 10178 4326 10190 4378
rect 10242 4326 10254 4378
rect 10306 4326 10318 4378
rect 10370 4326 10764 4378
rect 1104 4304 10764 4326
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 7282 4264 7288 4276
rect 7239 4236 7288 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8159 4236 9996 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 5994 4196 6000 4208
rect 3476 4168 6000 4196
rect 3476 4156 3482 4168
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 3436 4100 4169 4128
rect 3436 4069 3464 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 5534 4128 5540 4140
rect 4663 4100 5540 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 3970 4060 3976 4072
rect 3743 4032 3976 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4172 4060 4200 4091
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 7466 4088 7472 4140
rect 7524 4088 7530 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 4430 4060 4436 4072
rect 4172 4032 4436 4060
rect 4065 4023 4123 4029
rect 4080 3992 4108 4023
rect 4430 4020 4436 4032
rect 4488 4060 4494 4072
rect 4525 4063 4583 4069
rect 4525 4060 4537 4063
rect 4488 4032 4537 4060
rect 4488 4020 4494 4032
rect 4525 4029 4537 4032
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4060 5043 4063
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5031 4032 5181 4060
rect 5031 4029 5043 4032
rect 4985 4023 5043 4029
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 7576 4060 7604 4091
rect 5169 4023 5227 4029
rect 7484 4032 7604 4060
rect 7653 4063 7711 4069
rect 4890 3992 4896 4004
rect 2746 3964 3832 3992
rect 4080 3964 4896 3992
rect 2746 3936 2774 3964
rect 2682 3884 2688 3936
rect 2740 3896 2774 3936
rect 3804 3933 3832 3964
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 7484 3992 7512 4032
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 7834 4060 7840 4072
rect 7699 4032 7840 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 7944 3992 7972 4091
rect 8754 4088 8760 4140
rect 8812 4088 8818 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 9858 4128 9864 4140
rect 9815 4100 9864 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9968 4128 9996 4236
rect 10594 4128 10600 4140
rect 9968 4100 10600 4128
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8895 4063 8953 4069
rect 8895 4060 8907 4063
rect 8628 4032 8907 4060
rect 8628 4020 8634 4032
rect 8895 4029 8907 4032
rect 8941 4029 8953 4063
rect 8895 4023 8953 4029
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9950 4020 9956 4072
rect 10008 4020 10014 4072
rect 7432 3964 7512 3992
rect 7668 3964 7972 3992
rect 7432 3952 7438 3964
rect 3789 3927 3847 3933
rect 2740 3884 2746 3896
rect 3789 3893 3801 3927
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5776 3896 5825 3924
rect 5776 3884 5782 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7668 3924 7696 3964
rect 7524 3896 7696 3924
rect 7524 3884 7530 3896
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 7944 3924 7972 3964
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 8938 3924 8944 3936
rect 7944 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3924 9002 3936
rect 9324 3924 9352 3955
rect 8996 3896 9352 3924
rect 8996 3884 9002 3896
rect 1104 3834 10764 3856
rect 1104 3782 2157 3834
rect 2209 3782 2221 3834
rect 2273 3782 2285 3834
rect 2337 3782 2349 3834
rect 2401 3782 2413 3834
rect 2465 3782 4572 3834
rect 4624 3782 4636 3834
rect 4688 3782 4700 3834
rect 4752 3782 4764 3834
rect 4816 3782 4828 3834
rect 4880 3782 6987 3834
rect 7039 3782 7051 3834
rect 7103 3782 7115 3834
rect 7167 3782 7179 3834
rect 7231 3782 7243 3834
rect 7295 3782 9402 3834
rect 9454 3782 9466 3834
rect 9518 3782 9530 3834
rect 9582 3782 9594 3834
rect 9646 3782 9658 3834
rect 9710 3782 10764 3834
rect 1104 3760 10764 3782
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3384 3692 4537 3720
rect 3384 3680 3390 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 5524 3723 5582 3729
rect 5524 3689 5536 3723
rect 5570 3720 5582 3723
rect 5718 3720 5724 3732
rect 5570 3692 5724 3720
rect 5570 3689 5582 3692
rect 5524 3683 5582 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7466 3720 7472 3732
rect 7055 3692 7472 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 8481 3723 8539 3729
rect 7800 3692 8248 3720
rect 7800 3680 7806 3692
rect 8220 3664 8248 3692
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8570 3720 8576 3732
rect 8527 3692 8576 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10410 3720 10416 3732
rect 10008 3692 10416 3720
rect 10008 3680 10014 3692
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 8260 3624 8677 3652
rect 8260 3612 8266 3624
rect 8665 3621 8677 3624
rect 8711 3621 8723 3655
rect 8665 3615 8723 3621
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1946 3584 1952 3596
rect 1627 3556 1952 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1946 3544 1952 3556
rect 2004 3584 2010 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 2004 3556 5273 3584
rect 2004 3544 2010 3556
rect 3712 3528 3740 3556
rect 5261 3553 5273 3556
rect 5307 3584 5319 3587
rect 5626 3584 5632 3596
rect 5307 3556 5632 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5626 3544 5632 3556
rect 5684 3584 5690 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 5684 3556 7113 3584
rect 5684 3544 5690 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 8478 3584 8484 3596
rect 7101 3547 7159 3553
rect 8128 3556 8484 3584
rect 3418 3516 3424 3528
rect 2990 3488 3424 3516
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3694 3476 3700 3528
rect 3752 3476 3758 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 7116 3516 7144 3547
rect 8128 3516 8156 3556
rect 8478 3544 8484 3556
rect 8536 3584 8542 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8536 3556 9045 3584
rect 8536 3544 8542 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 7116 3488 8156 3516
rect 1854 3408 1860 3460
rect 1912 3408 1918 3460
rect 4356 3448 4384 3479
rect 3344 3420 4384 3448
rect 3344 3389 3372 3420
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3349 3387 3383
rect 3329 3343 3387 3349
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 5184 3380 5212 3479
rect 5994 3408 6000 3460
rect 6052 3408 6058 3460
rect 5626 3380 5632 3392
rect 5184 3352 5632 3380
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 7116 3380 7144 3488
rect 8754 3476 8760 3528
rect 8812 3476 8818 3528
rect 7368 3451 7426 3457
rect 7368 3417 7380 3451
rect 7414 3448 7426 3451
rect 7558 3448 7564 3460
rect 7414 3420 7564 3448
rect 7414 3417 7426 3420
rect 7368 3411 7426 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 7282 3380 7288 3392
rect 7116 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8772 3380 8800 3476
rect 9300 3451 9358 3457
rect 9300 3417 9312 3451
rect 9346 3448 9358 3451
rect 9858 3448 9864 3460
rect 9346 3420 9864 3448
rect 9346 3417 9358 3420
rect 9300 3411 9358 3417
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 7524 3352 8800 3380
rect 7524 3340 7530 3352
rect 1104 3290 10764 3312
rect 1104 3238 2817 3290
rect 2869 3238 2881 3290
rect 2933 3238 2945 3290
rect 2997 3238 3009 3290
rect 3061 3238 3073 3290
rect 3125 3238 5232 3290
rect 5284 3238 5296 3290
rect 5348 3238 5360 3290
rect 5412 3238 5424 3290
rect 5476 3238 5488 3290
rect 5540 3238 7647 3290
rect 7699 3238 7711 3290
rect 7763 3238 7775 3290
rect 7827 3238 7839 3290
rect 7891 3238 7903 3290
rect 7955 3238 10062 3290
rect 10114 3238 10126 3290
rect 10178 3238 10190 3290
rect 10242 3238 10254 3290
rect 10306 3238 10318 3290
rect 10370 3238 10764 3290
rect 1104 3216 10764 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 2409 3179 2467 3185
rect 2409 3176 2421 3179
rect 1912 3148 2421 3176
rect 1912 3136 1918 3148
rect 2409 3145 2421 3148
rect 2455 3145 2467 3179
rect 2409 3139 2467 3145
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 8294 3176 8300 3188
rect 7208 3148 8300 3176
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3804 3040 3832 3136
rect 6178 3068 6184 3120
rect 6236 3068 6242 3120
rect 7208 3049 7236 3148
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9030 3136 9036 3188
rect 9088 3136 9094 3188
rect 9858 3136 9864 3188
rect 9916 3136 9922 3188
rect 10229 3179 10287 3185
rect 10229 3145 10241 3179
rect 10275 3176 10287 3179
rect 10686 3176 10692 3188
rect 10275 3148 10692 3176
rect 10275 3145 10287 3148
rect 10229 3139 10287 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 7561 3111 7619 3117
rect 7561 3077 7573 3111
rect 7607 3108 7619 3111
rect 7607 3080 9260 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 3559 3012 3832 3040
rect 7101 3043 7159 3049
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3142 2972 3148 2984
rect 3007 2944 3148 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 5626 2972 5632 2984
rect 3651 2944 5632 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4062 2904 4068 2916
rect 3476 2876 4068 2904
rect 3476 2864 3482 2876
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 3752 2808 4721 2836
rect 3752 2796 3758 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 7116 2836 7144 3003
rect 7300 2972 7328 3068
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7466 3040 7472 3052
rect 7423 3012 7472 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7926 3049 7932 3052
rect 7920 3003 7932 3049
rect 7926 3000 7932 3003
rect 7984 3000 7990 3052
rect 9232 3049 9260 3080
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3040 10471 3043
rect 10888 3040 10916 3136
rect 10459 3012 10916 3040
rect 10459 3009 10471 3012
rect 10413 3003 10471 3009
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7300 2944 7665 2972
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 7374 2904 7380 2916
rect 7331 2876 7380 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 9766 2836 9772 2848
rect 7116 2808 9772 2836
rect 4709 2799 4767 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 1104 2746 10764 2768
rect 1104 2694 2157 2746
rect 2209 2694 2221 2746
rect 2273 2694 2285 2746
rect 2337 2694 2349 2746
rect 2401 2694 2413 2746
rect 2465 2694 4572 2746
rect 4624 2694 4636 2746
rect 4688 2694 4700 2746
rect 4752 2694 4764 2746
rect 4816 2694 4828 2746
rect 4880 2694 6987 2746
rect 7039 2694 7051 2746
rect 7103 2694 7115 2746
rect 7167 2694 7179 2746
rect 7231 2694 7243 2746
rect 7295 2694 9402 2746
rect 9454 2694 9466 2746
rect 9518 2694 9530 2746
rect 9582 2694 9594 2746
rect 9646 2694 9658 2746
rect 9710 2694 10764 2746
rect 1104 2672 10764 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 3234 2632 3240 2644
rect 3099 2604 3240 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7984 2604 8033 2632
rect 7984 2592 7990 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8021 2595 8079 2601
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3752 2468 3801 2496
rect 3752 2456 3758 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 7392 2496 7420 2592
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 8389 2567 8447 2573
rect 8389 2564 8401 2567
rect 8352 2536 8401 2564
rect 8352 2524 8358 2536
rect 8389 2533 8401 2536
rect 8435 2533 8447 2567
rect 8389 2527 8447 2533
rect 7392 2468 8340 2496
rect 3789 2459 3847 2465
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 4028 2332 4077 2360
rect 4028 2320 4034 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 4065 2323 4123 2329
rect 4338 2320 4344 2372
rect 4396 2360 4402 2372
rect 7760 2360 7788 2391
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8312 2437 8340 2468
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9088 2468 9505 2496
rect 9088 2456 9094 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 10410 2456 10416 2508
rect 10468 2456 10474 2508
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8527 2400 8953 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 8754 2360 8760 2372
rect 4396 2332 4554 2360
rect 7760 2332 8760 2360
rect 4396 2320 4402 2332
rect 8754 2320 8760 2332
rect 8812 2320 8818 2372
rect 7929 2295 7987 2301
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8662 2292 8668 2304
rect 7975 2264 8668 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 1104 2202 10764 2224
rect 1104 2150 2817 2202
rect 2869 2150 2881 2202
rect 2933 2150 2945 2202
rect 2997 2150 3009 2202
rect 3061 2150 3073 2202
rect 3125 2150 5232 2202
rect 5284 2150 5296 2202
rect 5348 2150 5360 2202
rect 5412 2150 5424 2202
rect 5476 2150 5488 2202
rect 5540 2150 7647 2202
rect 7699 2150 7711 2202
rect 7763 2150 7775 2202
rect 7827 2150 7839 2202
rect 7891 2150 7903 2202
rect 7955 2150 10062 2202
rect 10114 2150 10126 2202
rect 10178 2150 10190 2202
rect 10242 2150 10254 2202
rect 10306 2150 10318 2202
rect 10370 2150 10764 2202
rect 1104 2128 10764 2150
<< via1 >>
rect 2157 11398 2209 11450
rect 2221 11398 2273 11450
rect 2285 11398 2337 11450
rect 2349 11398 2401 11450
rect 2413 11398 2465 11450
rect 4572 11398 4624 11450
rect 4636 11398 4688 11450
rect 4700 11398 4752 11450
rect 4764 11398 4816 11450
rect 4828 11398 4880 11450
rect 6987 11398 7039 11450
rect 7051 11398 7103 11450
rect 7115 11398 7167 11450
rect 7179 11398 7231 11450
rect 7243 11398 7295 11450
rect 9402 11398 9454 11450
rect 9466 11398 9518 11450
rect 9530 11398 9582 11450
rect 9594 11398 9646 11450
rect 9658 11398 9710 11450
rect 2964 11296 3016 11348
rect 8944 11296 8996 11348
rect 4252 11092 4304 11144
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 3148 11024 3200 11033
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 7380 11024 7432 11076
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 3332 10956 3384 11008
rect 8208 10956 8260 11008
rect 2817 10854 2869 10906
rect 2881 10854 2933 10906
rect 2945 10854 2997 10906
rect 3009 10854 3061 10906
rect 3073 10854 3125 10906
rect 5232 10854 5284 10906
rect 5296 10854 5348 10906
rect 5360 10854 5412 10906
rect 5424 10854 5476 10906
rect 5488 10854 5540 10906
rect 7647 10854 7699 10906
rect 7711 10854 7763 10906
rect 7775 10854 7827 10906
rect 7839 10854 7891 10906
rect 7903 10854 7955 10906
rect 10062 10854 10114 10906
rect 10126 10854 10178 10906
rect 10190 10854 10242 10906
rect 10254 10854 10306 10906
rect 10318 10854 10370 10906
rect 3148 10752 3200 10804
rect 940 10616 992 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 8116 10752 8168 10804
rect 9128 10752 9180 10804
rect 8392 10684 8444 10736
rect 4436 10548 4488 10600
rect 6920 10616 6972 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7748 10616 7800 10668
rect 3608 10480 3660 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 3700 10412 3752 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5816 10548 5868 10600
rect 7656 10548 7708 10600
rect 5632 10412 5684 10464
rect 5724 10412 5776 10464
rect 7564 10412 7616 10464
rect 8668 10616 8720 10668
rect 10876 10480 10928 10532
rect 9220 10412 9272 10464
rect 2157 10310 2209 10362
rect 2221 10310 2273 10362
rect 2285 10310 2337 10362
rect 2349 10310 2401 10362
rect 2413 10310 2465 10362
rect 4572 10310 4624 10362
rect 4636 10310 4688 10362
rect 4700 10310 4752 10362
rect 4764 10310 4816 10362
rect 4828 10310 4880 10362
rect 6987 10310 7039 10362
rect 7051 10310 7103 10362
rect 7115 10310 7167 10362
rect 7179 10310 7231 10362
rect 7243 10310 7295 10362
rect 9402 10310 9454 10362
rect 9466 10310 9518 10362
rect 9530 10310 9582 10362
rect 9594 10310 9646 10362
rect 9658 10310 9710 10362
rect 1584 10208 1636 10260
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3424 10208 3476 10260
rect 5724 10208 5776 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 3608 10004 3660 10056
rect 5632 10072 5684 10124
rect 7748 10072 7800 10124
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 3700 9936 3752 9988
rect 4712 9936 4764 9988
rect 3884 9868 3936 9920
rect 6828 10004 6880 10056
rect 6552 9979 6604 9988
rect 6552 9945 6586 9979
rect 6586 9945 6604 9979
rect 6552 9936 6604 9945
rect 7104 9936 7156 9988
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8484 10072 8536 10124
rect 9220 10072 9272 10124
rect 10692 10208 10744 10260
rect 7380 9868 7432 9920
rect 9496 9868 9548 9920
rect 2817 9766 2869 9818
rect 2881 9766 2933 9818
rect 2945 9766 2997 9818
rect 3009 9766 3061 9818
rect 3073 9766 3125 9818
rect 5232 9766 5284 9818
rect 5296 9766 5348 9818
rect 5360 9766 5412 9818
rect 5424 9766 5476 9818
rect 5488 9766 5540 9818
rect 7647 9766 7699 9818
rect 7711 9766 7763 9818
rect 7775 9766 7827 9818
rect 7839 9766 7891 9818
rect 7903 9766 7955 9818
rect 10062 9766 10114 9818
rect 10126 9766 10178 9818
rect 10190 9766 10242 9818
rect 10254 9766 10306 9818
rect 10318 9766 10370 9818
rect 2688 9664 2740 9716
rect 3608 9664 3660 9716
rect 4712 9664 4764 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 6644 9664 6696 9716
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 8484 9664 8536 9716
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 5724 9528 5776 9580
rect 7104 9528 7156 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7472 9528 7524 9580
rect 9496 9596 9548 9648
rect 4436 9460 4488 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 6920 9460 6972 9512
rect 8116 9460 8168 9512
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 4252 9392 4304 9444
rect 5448 9392 5500 9444
rect 6000 9324 6052 9376
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 8208 9324 8260 9376
rect 2157 9222 2209 9274
rect 2221 9222 2273 9274
rect 2285 9222 2337 9274
rect 2349 9222 2401 9274
rect 2413 9222 2465 9274
rect 4572 9222 4624 9274
rect 4636 9222 4688 9274
rect 4700 9222 4752 9274
rect 4764 9222 4816 9274
rect 4828 9222 4880 9274
rect 6987 9222 7039 9274
rect 7051 9222 7103 9274
rect 7115 9222 7167 9274
rect 7179 9222 7231 9274
rect 7243 9222 7295 9274
rect 9402 9222 9454 9274
rect 9466 9222 9518 9274
rect 9530 9222 9582 9274
rect 9594 9222 9646 9274
rect 9658 9222 9710 9274
rect 3608 9120 3660 9172
rect 4436 9120 4488 9172
rect 5080 9120 5132 9172
rect 5724 9120 5776 9172
rect 5448 8916 5500 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6644 9052 6696 9104
rect 5632 8848 5684 8900
rect 7380 8848 7432 8900
rect 6920 8780 6972 8832
rect 8024 8891 8076 8900
rect 8024 8857 8033 8891
rect 8033 8857 8067 8891
rect 8067 8857 8076 8891
rect 8024 8848 8076 8857
rect 9864 8848 9916 8900
rect 8116 8780 8168 8832
rect 9220 8780 9272 8832
rect 2817 8678 2869 8730
rect 2881 8678 2933 8730
rect 2945 8678 2997 8730
rect 3009 8678 3061 8730
rect 3073 8678 3125 8730
rect 5232 8678 5284 8730
rect 5296 8678 5348 8730
rect 5360 8678 5412 8730
rect 5424 8678 5476 8730
rect 5488 8678 5540 8730
rect 7647 8678 7699 8730
rect 7711 8678 7763 8730
rect 7775 8678 7827 8730
rect 7839 8678 7891 8730
rect 7903 8678 7955 8730
rect 10062 8678 10114 8730
rect 10126 8678 10178 8730
rect 10190 8678 10242 8730
rect 10254 8678 10306 8730
rect 10318 8678 10370 8730
rect 6736 8576 6788 8628
rect 8392 8576 8444 8628
rect 9036 8576 9088 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 3332 8440 3384 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 6828 8508 6880 8560
rect 6920 8440 6972 8492
rect 8024 8440 8076 8492
rect 8208 8483 8260 8492
rect 8208 8449 8242 8483
rect 8242 8449 8260 8483
rect 8208 8440 8260 8449
rect 3976 8304 4028 8356
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 6276 8236 6328 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 2157 8134 2209 8186
rect 2221 8134 2273 8186
rect 2285 8134 2337 8186
rect 2349 8134 2401 8186
rect 2413 8134 2465 8186
rect 4572 8134 4624 8186
rect 4636 8134 4688 8186
rect 4700 8134 4752 8186
rect 4764 8134 4816 8186
rect 4828 8134 4880 8186
rect 6987 8134 7039 8186
rect 7051 8134 7103 8186
rect 7115 8134 7167 8186
rect 7179 8134 7231 8186
rect 7243 8134 7295 8186
rect 9402 8134 9454 8186
rect 9466 8134 9518 8186
rect 9530 8134 9582 8186
rect 9594 8134 9646 8186
rect 9658 8134 9710 8186
rect 1860 8032 1912 8084
rect 6828 8032 6880 8084
rect 6092 7964 6144 8016
rect 7472 8032 7524 8084
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 3148 7896 3200 7948
rect 3884 7896 3936 7948
rect 9128 7896 9180 7948
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 6276 7828 6328 7880
rect 7564 7828 7616 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 10600 7896 10652 7948
rect 3608 7760 3660 7812
rect 6184 7760 6236 7812
rect 8024 7692 8076 7744
rect 8300 7692 8352 7744
rect 9772 7692 9824 7744
rect 9864 7692 9916 7744
rect 9956 7692 10008 7744
rect 10416 7692 10468 7744
rect 2817 7590 2869 7642
rect 2881 7590 2933 7642
rect 2945 7590 2997 7642
rect 3009 7590 3061 7642
rect 3073 7590 3125 7642
rect 5232 7590 5284 7642
rect 5296 7590 5348 7642
rect 5360 7590 5412 7642
rect 5424 7590 5476 7642
rect 5488 7590 5540 7642
rect 7647 7590 7699 7642
rect 7711 7590 7763 7642
rect 7775 7590 7827 7642
rect 7839 7590 7891 7642
rect 7903 7590 7955 7642
rect 10062 7590 10114 7642
rect 10126 7590 10178 7642
rect 10190 7590 10242 7642
rect 10254 7590 10306 7642
rect 10318 7590 10370 7642
rect 1584 7352 1636 7404
rect 2688 7488 2740 7540
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 3332 7352 3384 7404
rect 6828 7488 6880 7540
rect 7564 7488 7616 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 8576 7488 8628 7540
rect 9220 7488 9272 7540
rect 3148 7284 3200 7336
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 5632 7352 5684 7404
rect 6276 7352 6328 7404
rect 8116 7420 8168 7472
rect 6092 7284 6144 7336
rect 8392 7352 8444 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 10416 7352 10468 7404
rect 8576 7284 8628 7336
rect 9128 7284 9180 7336
rect 9864 7284 9916 7336
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10508 7148 10560 7200
rect 2157 7046 2209 7098
rect 2221 7046 2273 7098
rect 2285 7046 2337 7098
rect 2349 7046 2401 7098
rect 2413 7046 2465 7098
rect 4572 7046 4624 7098
rect 4636 7046 4688 7098
rect 4700 7046 4752 7098
rect 4764 7046 4816 7098
rect 4828 7046 4880 7098
rect 6987 7046 7039 7098
rect 7051 7046 7103 7098
rect 7115 7046 7167 7098
rect 7179 7046 7231 7098
rect 7243 7046 7295 7098
rect 9402 7046 9454 7098
rect 9466 7046 9518 7098
rect 9530 7046 9582 7098
rect 9594 7046 9646 7098
rect 9658 7046 9710 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 3608 6944 3660 6996
rect 8576 6944 8628 6996
rect 1860 6808 1912 6860
rect 3148 6808 3200 6860
rect 3332 6808 3384 6860
rect 5540 6808 5592 6860
rect 10324 6876 10376 6928
rect 9864 6808 9916 6860
rect 3424 6740 3476 6792
rect 4160 6672 4212 6724
rect 7472 6672 7524 6724
rect 3148 6604 3200 6656
rect 6184 6604 6236 6656
rect 8484 6604 8536 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 2817 6502 2869 6554
rect 2881 6502 2933 6554
rect 2945 6502 2997 6554
rect 3009 6502 3061 6554
rect 3073 6502 3125 6554
rect 5232 6502 5284 6554
rect 5296 6502 5348 6554
rect 5360 6502 5412 6554
rect 5424 6502 5476 6554
rect 5488 6502 5540 6554
rect 7647 6502 7699 6554
rect 7711 6502 7763 6554
rect 7775 6502 7827 6554
rect 7839 6502 7891 6554
rect 7903 6502 7955 6554
rect 10062 6502 10114 6554
rect 10126 6502 10178 6554
rect 10190 6502 10242 6554
rect 10254 6502 10306 6554
rect 10318 6502 10370 6554
rect 7472 6400 7524 6452
rect 8024 6400 8076 6452
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4896 6264 4948 6316
rect 5632 6264 5684 6316
rect 9680 6400 9732 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 8392 6264 8444 6316
rect 3332 6196 3384 6248
rect 3608 6196 3660 6248
rect 5632 6060 5684 6112
rect 5816 6060 5868 6112
rect 6000 6060 6052 6112
rect 8484 6060 8536 6112
rect 2157 5958 2209 6010
rect 2221 5958 2273 6010
rect 2285 5958 2337 6010
rect 2349 5958 2401 6010
rect 2413 5958 2465 6010
rect 4572 5958 4624 6010
rect 4636 5958 4688 6010
rect 4700 5958 4752 6010
rect 4764 5958 4816 6010
rect 4828 5958 4880 6010
rect 6987 5958 7039 6010
rect 7051 5958 7103 6010
rect 7115 5958 7167 6010
rect 7179 5958 7231 6010
rect 7243 5958 7295 6010
rect 9402 5958 9454 6010
rect 9466 5958 9518 6010
rect 9530 5958 9582 6010
rect 9594 5958 9646 6010
rect 9658 5958 9710 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 8116 5856 8168 5908
rect 9956 5856 10008 5908
rect 3148 5720 3200 5772
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 3056 5652 3108 5704
rect 3976 5652 4028 5704
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10508 5584 10560 5636
rect 2228 5516 2280 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 4896 5516 4948 5568
rect 5632 5516 5684 5568
rect 6000 5516 6052 5568
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 8944 5516 8996 5568
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 9864 5516 9916 5568
rect 2817 5414 2869 5466
rect 2881 5414 2933 5466
rect 2945 5414 2997 5466
rect 3009 5414 3061 5466
rect 3073 5414 3125 5466
rect 5232 5414 5284 5466
rect 5296 5414 5348 5466
rect 5360 5414 5412 5466
rect 5424 5414 5476 5466
rect 5488 5414 5540 5466
rect 7647 5414 7699 5466
rect 7711 5414 7763 5466
rect 7775 5414 7827 5466
rect 7839 5414 7891 5466
rect 7903 5414 7955 5466
rect 10062 5414 10114 5466
rect 10126 5414 10178 5466
rect 10190 5414 10242 5466
rect 10254 5414 10306 5466
rect 10318 5414 10370 5466
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 4712 5312 4764 5364
rect 6000 5312 6052 5364
rect 5724 5244 5776 5296
rect 9220 5244 9272 5296
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 2688 5108 2740 5160
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 3424 4972 3476 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 5632 4972 5684 5024
rect 8760 4972 8812 5024
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 2157 4870 2209 4922
rect 2221 4870 2273 4922
rect 2285 4870 2337 4922
rect 2349 4870 2401 4922
rect 2413 4870 2465 4922
rect 4572 4870 4624 4922
rect 4636 4870 4688 4922
rect 4700 4870 4752 4922
rect 4764 4870 4816 4922
rect 4828 4870 4880 4922
rect 6987 4870 7039 4922
rect 7051 4870 7103 4922
rect 7115 4870 7167 4922
rect 7179 4870 7231 4922
rect 7243 4870 7295 4922
rect 9402 4870 9454 4922
rect 9466 4870 9518 4922
rect 9530 4870 9582 4922
rect 9594 4870 9646 4922
rect 9658 4870 9710 4922
rect 3700 4768 3752 4820
rect 8116 4768 8168 4820
rect 9772 4768 9824 4820
rect 7380 4700 7432 4752
rect 9864 4632 9916 4684
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 7472 4564 7524 4616
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 8760 4564 8812 4616
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 4436 4428 4488 4480
rect 7564 4428 7616 4480
rect 2817 4326 2869 4378
rect 2881 4326 2933 4378
rect 2945 4326 2997 4378
rect 3009 4326 3061 4378
rect 3073 4326 3125 4378
rect 5232 4326 5284 4378
rect 5296 4326 5348 4378
rect 5360 4326 5412 4378
rect 5424 4326 5476 4378
rect 5488 4326 5540 4378
rect 7647 4326 7699 4378
rect 7711 4326 7763 4378
rect 7775 4326 7827 4378
rect 7839 4326 7891 4378
rect 7903 4326 7955 4378
rect 10062 4326 10114 4378
rect 10126 4326 10178 4378
rect 10190 4326 10242 4378
rect 10254 4326 10306 4378
rect 10318 4326 10370 4378
rect 7288 4224 7340 4276
rect 3424 4156 3476 4208
rect 6000 4156 6052 4208
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3976 4020 4028 4072
rect 5540 4088 5592 4140
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 4436 4020 4488 4072
rect 2688 3884 2740 3936
rect 4896 3952 4948 4004
rect 7380 3952 7432 4004
rect 7840 4020 7892 4072
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9864 4088 9916 4140
rect 10600 4088 10652 4140
rect 8576 4020 8628 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 5724 3884 5776 3936
rect 7472 3884 7524 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8944 3884 8996 3936
rect 2157 3782 2209 3834
rect 2221 3782 2273 3834
rect 2285 3782 2337 3834
rect 2349 3782 2401 3834
rect 2413 3782 2465 3834
rect 4572 3782 4624 3834
rect 4636 3782 4688 3834
rect 4700 3782 4752 3834
rect 4764 3782 4816 3834
rect 4828 3782 4880 3834
rect 6987 3782 7039 3834
rect 7051 3782 7103 3834
rect 7115 3782 7167 3834
rect 7179 3782 7231 3834
rect 7243 3782 7295 3834
rect 9402 3782 9454 3834
rect 9466 3782 9518 3834
rect 9530 3782 9582 3834
rect 9594 3782 9646 3834
rect 9658 3782 9710 3834
rect 3332 3680 3384 3732
rect 5724 3680 5776 3732
rect 7472 3680 7524 3732
rect 7748 3680 7800 3732
rect 8576 3680 8628 3732
rect 9956 3680 10008 3732
rect 10416 3723 10468 3732
rect 10416 3689 10425 3723
rect 10425 3689 10459 3723
rect 10459 3689 10468 3723
rect 10416 3680 10468 3689
rect 8208 3612 8260 3664
rect 1952 3544 2004 3596
rect 5632 3544 5684 3596
rect 3424 3476 3476 3528
rect 3700 3476 3752 3528
rect 8484 3544 8536 3596
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 6000 3408 6052 3460
rect 5632 3340 5684 3392
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 7564 3408 7616 3460
rect 7288 3340 7340 3392
rect 7472 3340 7524 3392
rect 9864 3408 9916 3460
rect 2817 3238 2869 3290
rect 2881 3238 2933 3290
rect 2945 3238 2997 3290
rect 3009 3238 3061 3290
rect 3073 3238 3125 3290
rect 5232 3238 5284 3290
rect 5296 3238 5348 3290
rect 5360 3238 5412 3290
rect 5424 3238 5476 3290
rect 5488 3238 5540 3290
rect 7647 3238 7699 3290
rect 7711 3238 7763 3290
rect 7775 3238 7827 3290
rect 7839 3238 7891 3290
rect 7903 3238 7955 3290
rect 10062 3238 10114 3290
rect 10126 3238 10178 3290
rect 10190 3238 10242 3290
rect 10254 3238 10306 3290
rect 10318 3238 10370 3290
rect 1860 3136 1912 3188
rect 3792 3136 3844 3188
rect 6184 3111 6236 3120
rect 6184 3077 6193 3111
rect 6193 3077 6227 3111
rect 6227 3077 6236 3111
rect 6184 3068 6236 3077
rect 8300 3136 8352 3188
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10692 3136 10744 3188
rect 10876 3136 10928 3188
rect 7288 3068 7340 3120
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 5632 2932 5684 2984
rect 3424 2864 3476 2916
rect 4068 2864 4120 2916
rect 3700 2796 3752 2848
rect 7472 3000 7524 3052
rect 7932 3043 7984 3052
rect 7932 3009 7966 3043
rect 7966 3009 7984 3043
rect 7932 3000 7984 3009
rect 7380 2864 7432 2916
rect 9772 2796 9824 2848
rect 2157 2694 2209 2746
rect 2221 2694 2273 2746
rect 2285 2694 2337 2746
rect 2349 2694 2401 2746
rect 2413 2694 2465 2746
rect 4572 2694 4624 2746
rect 4636 2694 4688 2746
rect 4700 2694 4752 2746
rect 4764 2694 4816 2746
rect 4828 2694 4880 2746
rect 6987 2694 7039 2746
rect 7051 2694 7103 2746
rect 7115 2694 7167 2746
rect 7179 2694 7231 2746
rect 7243 2694 7295 2746
rect 9402 2694 9454 2746
rect 9466 2694 9518 2746
rect 9530 2694 9582 2746
rect 9594 2694 9646 2746
rect 9658 2694 9710 2746
rect 3240 2592 3292 2644
rect 5632 2592 5684 2644
rect 7380 2592 7432 2644
rect 7932 2592 7984 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 3700 2456 3752 2508
rect 8300 2524 8352 2576
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3976 2320 4028 2372
rect 4344 2320 4396 2372
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 9036 2456 9088 2508
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 8760 2320 8812 2372
rect 8668 2252 8720 2304
rect 2817 2150 2869 2202
rect 2881 2150 2933 2202
rect 2945 2150 2997 2202
rect 3009 2150 3061 2202
rect 3073 2150 3125 2202
rect 5232 2150 5284 2202
rect 5296 2150 5348 2202
rect 5360 2150 5412 2202
rect 5424 2150 5476 2202
rect 5488 2150 5540 2202
rect 7647 2150 7699 2202
rect 7711 2150 7763 2202
rect 7775 2150 7827 2202
rect 7839 2150 7891 2202
rect 7903 2150 7955 2202
rect 10062 2150 10114 2202
rect 10126 2150 10178 2202
rect 10190 2150 10242 2202
rect 10254 2150 10306 2202
rect 10318 2150 10370 2202
<< metal2 >>
rect 2962 13298 3018 14098
rect 8942 13298 8998 14098
rect 2157 11452 2465 11461
rect 2157 11450 2163 11452
rect 2219 11450 2243 11452
rect 2299 11450 2323 11452
rect 2379 11450 2403 11452
rect 2459 11450 2465 11452
rect 2219 11398 2221 11450
rect 2401 11398 2403 11450
rect 2157 11396 2163 11398
rect 2219 11396 2243 11398
rect 2299 11396 2323 11398
rect 2379 11396 2403 11398
rect 2459 11396 2465 11398
rect 2157 11387 2465 11396
rect 2976 11354 3004 13298
rect 4572 11452 4880 11461
rect 4572 11450 4578 11452
rect 4634 11450 4658 11452
rect 4714 11450 4738 11452
rect 4794 11450 4818 11452
rect 4874 11450 4880 11452
rect 4634 11398 4636 11450
rect 4816 11398 4818 11450
rect 4572 11396 4578 11398
rect 4634 11396 4658 11398
rect 4714 11396 4738 11398
rect 4794 11396 4818 11398
rect 4874 11396 4880 11398
rect 4572 11387 4880 11396
rect 6987 11452 7295 11461
rect 6987 11450 6993 11452
rect 7049 11450 7073 11452
rect 7129 11450 7153 11452
rect 7209 11450 7233 11452
rect 7289 11450 7295 11452
rect 7049 11398 7051 11450
rect 7231 11398 7233 11450
rect 6987 11396 6993 11398
rect 7049 11396 7073 11398
rect 7129 11396 7153 11398
rect 7209 11396 7233 11398
rect 7289 11396 7295 11398
rect 6987 11387 7295 11396
rect 8956 11354 8984 13298
rect 9402 11452 9710 11461
rect 9402 11450 9408 11452
rect 9464 11450 9488 11452
rect 9544 11450 9568 11452
rect 9624 11450 9648 11452
rect 9704 11450 9710 11452
rect 9464 11398 9466 11450
rect 9646 11398 9648 11450
rect 9402 11396 9408 11398
rect 9464 11396 9488 11398
rect 9544 11396 9568 11398
rect 9624 11396 9648 11398
rect 9704 11396 9710 11398
rect 9402 11387 9710 11396
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 2817 10908 3125 10917
rect 2817 10906 2823 10908
rect 2879 10906 2903 10908
rect 2959 10906 2983 10908
rect 3039 10906 3063 10908
rect 3119 10906 3125 10908
rect 2879 10854 2881 10906
rect 3061 10854 3063 10906
rect 2817 10852 2823 10854
rect 2879 10852 2903 10854
rect 2959 10852 2983 10854
rect 3039 10852 3063 10854
rect 3119 10852 3125 10854
rect 2817 10843 3125 10852
rect 3160 10810 3188 11018
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 952 10441 980 10610
rect 1584 10464 1636 10470
rect 938 10432 994 10441
rect 1584 10406 1636 10412
rect 938 10367 994 10376
rect 1596 10266 1624 10406
rect 2157 10364 2465 10373
rect 2157 10362 2163 10364
rect 2219 10362 2243 10364
rect 2299 10362 2323 10364
rect 2379 10362 2403 10364
rect 2459 10362 2465 10364
rect 2219 10310 2221 10362
rect 2401 10310 2403 10362
rect 2157 10308 2163 10310
rect 2219 10308 2243 10310
rect 2299 10308 2323 10310
rect 2379 10308 2403 10310
rect 2459 10308 2465 10310
rect 2157 10299 2465 10308
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 3068 9908 3096 10610
rect 3344 10266 3372 10950
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 10266 3464 10610
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3620 10062 3648 10474
rect 4264 10470 4292 11086
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 5232 10908 5540 10917
rect 5232 10906 5238 10908
rect 5294 10906 5318 10908
rect 5374 10906 5398 10908
rect 5454 10906 5478 10908
rect 5534 10906 5540 10908
rect 5294 10854 5296 10906
rect 5476 10854 5478 10906
rect 5232 10852 5238 10854
rect 5294 10852 5318 10854
rect 5374 10852 5398 10854
rect 5454 10852 5478 10854
rect 5534 10852 5540 10854
rect 5232 10843 5540 10852
rect 6932 10674 6960 11018
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3068 9880 3280 9908
rect 2817 9820 3125 9829
rect 2817 9818 2823 9820
rect 2879 9818 2903 9820
rect 2959 9818 2983 9820
rect 3039 9818 3063 9820
rect 3119 9818 3125 9820
rect 2879 9766 2881 9818
rect 3061 9766 3063 9818
rect 2817 9764 2823 9766
rect 2879 9764 2903 9766
rect 2959 9764 2983 9766
rect 3039 9764 3063 9766
rect 3119 9764 3125 9766
rect 2817 9755 3125 9764
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2157 9276 2465 9285
rect 2157 9274 2163 9276
rect 2219 9274 2243 9276
rect 2299 9274 2323 9276
rect 2379 9274 2403 9276
rect 2459 9274 2465 9276
rect 2219 9222 2221 9274
rect 2401 9222 2403 9274
rect 2157 9220 2163 9222
rect 2219 9220 2243 9222
rect 2299 9220 2323 9222
rect 2379 9220 2403 9222
rect 2459 9220 2465 9222
rect 2157 9211 2465 9220
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 7410 1624 8434
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 8090 1900 8366
rect 2157 8188 2465 8197
rect 2157 8186 2163 8188
rect 2219 8186 2243 8188
rect 2299 8186 2323 8188
rect 2379 8186 2403 8188
rect 2459 8186 2465 8188
rect 2219 8134 2221 8186
rect 2401 8134 2403 8186
rect 2157 8132 2163 8134
rect 2219 8132 2243 8134
rect 2299 8132 2323 8134
rect 2379 8132 2403 8134
rect 2459 8132 2465 8134
rect 2157 8123 2465 8132
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2700 7546 2728 9658
rect 2817 8732 3125 8741
rect 2817 8730 2823 8732
rect 2879 8730 2903 8732
rect 2959 8730 2983 8732
rect 3039 8730 3063 8732
rect 3119 8730 3125 8732
rect 2879 8678 2881 8730
rect 3061 8678 3063 8730
rect 2817 8676 2823 8678
rect 2879 8676 2903 8678
rect 2959 8676 2983 8678
rect 3039 8676 3063 8678
rect 3119 8676 3125 8678
rect 2817 8667 3125 8676
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2817 7644 3125 7653
rect 2817 7642 2823 7644
rect 2879 7642 2903 7644
rect 2959 7642 2983 7644
rect 3039 7642 3063 7644
rect 3119 7642 3125 7644
rect 2879 7590 2881 7642
rect 3061 7590 3063 7642
rect 2817 7588 2823 7590
rect 2879 7588 2903 7590
rect 2959 7588 2983 7590
rect 3039 7588 3063 7590
rect 3119 7588 3125 7590
rect 2817 7579 3125 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 3160 7342 3188 7890
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 1964 7002 1992 7278
rect 2157 7100 2465 7109
rect 2157 7098 2163 7100
rect 2219 7098 2243 7100
rect 2299 7098 2323 7100
rect 2379 7098 2403 7100
rect 2459 7098 2465 7100
rect 2219 7046 2221 7098
rect 2401 7046 2403 7098
rect 2157 7044 2163 7046
rect 2219 7044 2243 7046
rect 2299 7044 2323 7046
rect 2379 7044 2403 7046
rect 2459 7044 2465 7046
rect 2157 7035 2465 7044
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 3160 6866 3188 7278
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 1872 5914 1900 6802
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2817 6556 3125 6565
rect 2817 6554 2823 6556
rect 2879 6554 2903 6556
rect 2959 6554 2983 6556
rect 3039 6554 3063 6556
rect 3119 6554 3125 6556
rect 2879 6502 2881 6554
rect 3061 6502 3063 6554
rect 2817 6500 2823 6502
rect 2879 6500 2903 6502
rect 2959 6500 2983 6502
rect 3039 6500 3063 6502
rect 3119 6500 3125 6502
rect 2817 6491 3125 6500
rect 3160 6338 3188 6598
rect 3068 6310 3188 6338
rect 2157 6012 2465 6021
rect 2157 6010 2163 6012
rect 2219 6010 2243 6012
rect 2299 6010 2323 6012
rect 2379 6010 2403 6012
rect 2459 6010 2465 6012
rect 2219 5958 2221 6010
rect 2401 5958 2403 6010
rect 2157 5956 2163 5958
rect 2219 5956 2243 5958
rect 2299 5956 2323 5958
rect 2379 5956 2403 5958
rect 2459 5956 2465 5958
rect 2157 5947 2465 5956
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 3068 5710 3096 6310
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 5166 2268 5510
rect 2817 5468 3125 5477
rect 2817 5466 2823 5468
rect 2879 5466 2903 5468
rect 2959 5466 2983 5468
rect 3039 5466 3063 5468
rect 3119 5466 3125 5468
rect 2879 5414 2881 5466
rect 3061 5414 3063 5466
rect 2817 5412 2823 5414
rect 2879 5412 2903 5414
rect 2959 5412 2983 5414
rect 3039 5412 3063 5414
rect 3119 5412 3125 5414
rect 2817 5403 3125 5412
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1964 3602 1992 5102
rect 2157 4924 2465 4933
rect 2157 4922 2163 4924
rect 2219 4922 2243 4924
rect 2299 4922 2323 4924
rect 2379 4922 2403 4924
rect 2459 4922 2465 4924
rect 2219 4870 2221 4922
rect 2401 4870 2403 4922
rect 2157 4868 2163 4870
rect 2219 4868 2243 4870
rect 2299 4868 2323 4870
rect 2379 4868 2403 4870
rect 2459 4868 2465 4870
rect 2157 4859 2465 4868
rect 2700 3942 2728 5102
rect 2817 4380 3125 4389
rect 2817 4378 2823 4380
rect 2879 4378 2903 4380
rect 2959 4378 2983 4380
rect 3039 4378 3063 4380
rect 3119 4378 3125 4380
rect 2879 4326 2881 4378
rect 3061 4326 3063 4378
rect 2817 4324 2823 4326
rect 2879 4324 2903 4326
rect 2959 4324 2983 4326
rect 3039 4324 3063 4326
rect 3119 4324 3125 4326
rect 2817 4315 3125 4324
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2157 3836 2465 3845
rect 2157 3834 2163 3836
rect 2219 3834 2243 3836
rect 2299 3834 2323 3836
rect 2379 3834 2403 3836
rect 2459 3834 2465 3836
rect 2219 3782 2221 3834
rect 2401 3782 2403 3834
rect 2157 3780 2163 3782
rect 2219 3780 2243 3782
rect 2299 3780 2323 3782
rect 2379 3780 2403 3782
rect 2459 3780 2465 3782
rect 2157 3771 2465 3780
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1872 3194 1900 3402
rect 2817 3292 3125 3301
rect 2817 3290 2823 3292
rect 2879 3290 2903 3292
rect 2959 3290 2983 3292
rect 3039 3290 3063 3292
rect 3119 3290 3125 3292
rect 2879 3238 2881 3290
rect 3061 3238 3063 3290
rect 2817 3236 2823 3238
rect 2879 3236 2903 3238
rect 2959 3236 2983 3238
rect 3039 3236 3063 3238
rect 3119 3236 3125 3238
rect 2817 3227 3125 3236
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 3160 2990 3188 5714
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2157 2748 2465 2757
rect 2157 2746 2163 2748
rect 2219 2746 2243 2748
rect 2299 2746 2323 2748
rect 2379 2746 2403 2748
rect 2459 2746 2465 2748
rect 2219 2694 2221 2746
rect 2401 2694 2403 2746
rect 2157 2692 2163 2694
rect 2219 2692 2243 2694
rect 2299 2692 2323 2694
rect 2379 2692 2403 2694
rect 2459 2692 2465 2694
rect 2157 2683 2465 2692
rect 3252 2650 3280 9880
rect 3620 9722 3648 9998
rect 3712 9994 3740 10406
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3896 9586 3924 9862
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 4264 9450 4292 10406
rect 4448 9518 4476 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 4572 10364 4880 10373
rect 4572 10362 4578 10364
rect 4634 10362 4658 10364
rect 4714 10362 4738 10364
rect 4794 10362 4818 10364
rect 4874 10362 4880 10364
rect 4634 10310 4636 10362
rect 4816 10310 4818 10362
rect 4572 10308 4578 10310
rect 4634 10308 4658 10310
rect 4714 10308 4738 10310
rect 4794 10308 4818 10310
rect 4874 10308 4880 10310
rect 4572 10299 4880 10308
rect 5644 10130 5672 10406
rect 5736 10266 5764 10406
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4724 9722 4752 9930
rect 5232 9820 5540 9829
rect 5232 9818 5238 9820
rect 5294 9818 5318 9820
rect 5374 9818 5398 9820
rect 5454 9818 5478 9820
rect 5534 9818 5540 9820
rect 5294 9766 5296 9818
rect 5476 9766 5478 9818
rect 5232 9764 5238 9766
rect 5294 9764 5318 9766
rect 5374 9764 5398 9766
rect 5454 9764 5478 9766
rect 5534 9764 5540 9766
rect 5232 9755 5540 9764
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 5736 9586 5764 10202
rect 5828 10062 5856 10542
rect 6932 10418 6960 10610
rect 6840 10390 6960 10418
rect 6840 10282 6868 10390
rect 6987 10364 7295 10373
rect 6987 10362 6993 10364
rect 7049 10362 7073 10364
rect 7129 10362 7153 10364
rect 7209 10362 7233 10364
rect 7289 10362 7295 10364
rect 7049 10310 7051 10362
rect 7231 10310 7233 10362
rect 6987 10308 6993 10310
rect 7049 10308 7073 10310
rect 7129 10308 7153 10310
rect 7209 10308 7233 10310
rect 7289 10308 7295 10310
rect 6987 10299 7295 10308
rect 6840 10254 6960 10282
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9722 6592 9930
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6644 9716 6696 9722
rect 6840 9674 6868 9998
rect 6644 9658 6696 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9178 3648 9318
rect 4448 9178 4476 9454
rect 4572 9276 4880 9285
rect 4572 9274 4578 9276
rect 4634 9274 4658 9276
rect 4714 9274 4738 9276
rect 4794 9274 4818 9276
rect 4874 9274 4880 9276
rect 4634 9222 4636 9274
rect 4816 9222 4818 9274
rect 4572 9220 4578 9222
rect 4634 9220 4658 9222
rect 4714 9220 4738 9222
rect 4794 9220 4818 9222
rect 4874 9220 4880 9222
rect 4572 9211 4880 9220
rect 5092 9178 5120 9454
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5460 8974 5488 9386
rect 5736 9178 5764 9522
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 6012 8974 6040 9318
rect 6656 9110 6684 9658
rect 6748 9646 6868 9674
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5232 8732 5540 8741
rect 5232 8730 5238 8732
rect 5294 8730 5318 8732
rect 5374 8730 5398 8732
rect 5454 8730 5478 8732
rect 5534 8730 5540 8732
rect 5294 8678 5296 8730
rect 5476 8678 5478 8730
rect 5232 8676 5238 8678
rect 5294 8676 5318 8678
rect 5374 8676 5398 8678
rect 5454 8676 5478 8678
rect 5534 8676 5540 8678
rect 5232 8667 5540 8676
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 7410 3372 8434
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7954 3924 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3436 7290 3464 7822
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3344 7262 3464 7290
rect 3344 6866 3372 7262
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 6254 3372 6802
rect 3436 6798 3464 7142
rect 3620 7002 3648 7754
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3620 6254 3648 6938
rect 3988 6322 4016 8298
rect 4572 8188 4880 8197
rect 4572 8186 4578 8188
rect 4634 8186 4658 8188
rect 4714 8186 4738 8188
rect 4794 8186 4818 8188
rect 4874 8186 4880 8188
rect 4634 8134 4636 8186
rect 4816 8134 4818 8186
rect 4572 8132 4578 8134
rect 4634 8132 4658 8134
rect 4714 8132 4738 8134
rect 4794 8132 4818 8134
rect 4874 8132 4880 8134
rect 4572 8123 4880 8132
rect 5232 7644 5540 7653
rect 5232 7642 5238 7644
rect 5294 7642 5318 7644
rect 5374 7642 5398 7644
rect 5454 7642 5478 7644
rect 5534 7642 5540 7644
rect 5294 7590 5296 7642
rect 5476 7590 5478 7642
rect 5232 7588 5238 7590
rect 5294 7588 5318 7590
rect 5374 7588 5398 7590
rect 5454 7588 5478 7590
rect 5534 7588 5540 7590
rect 5232 7579 5540 7588
rect 5644 7410 5672 8842
rect 6748 8634 6776 9646
rect 6932 9518 6960 10254
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9586 7144 9930
rect 7392 9926 7420 11018
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7647 10908 7955 10917
rect 7647 10906 7653 10908
rect 7709 10906 7733 10908
rect 7789 10906 7813 10908
rect 7869 10906 7893 10908
rect 7949 10906 7955 10908
rect 7709 10854 7711 10906
rect 7891 10854 7893 10906
rect 7647 10852 7653 10854
rect 7709 10852 7733 10854
rect 7789 10852 7813 10854
rect 7869 10852 7893 10854
rect 7949 10852 7955 10854
rect 7647 10843 7955 10852
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9586 7420 9862
rect 7484 9586 7512 10610
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 9722 7604 10406
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7760 10130 7788 10610
rect 8128 10198 8156 10746
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7647 9820 7955 9829
rect 7647 9818 7653 9820
rect 7709 9818 7733 9820
rect 7789 9818 7813 9820
rect 7869 9818 7893 9820
rect 7949 9818 7955 9820
rect 7709 9766 7711 9818
rect 7891 9766 7893 9818
rect 7647 9764 7653 9766
rect 7709 9764 7733 9766
rect 7789 9764 7813 9766
rect 7869 9764 7893 9766
rect 7949 9764 7955 9766
rect 7647 9755 7955 9764
rect 8128 9722 8156 10134
rect 8220 10062 8248 10950
rect 9140 10810 9168 11018
rect 10062 10908 10370 10917
rect 10062 10906 10068 10908
rect 10124 10906 10148 10908
rect 10204 10906 10228 10908
rect 10284 10906 10308 10908
rect 10364 10906 10370 10908
rect 10124 10854 10126 10906
rect 10306 10854 10308 10906
rect 10062 10852 10068 10854
rect 10124 10852 10148 10854
rect 10204 10852 10228 10854
rect 10284 10852 10308 10854
rect 10364 10852 10370 10854
rect 10062 10843 10370 10852
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8404 10266 8432 10678
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 9330 6960 9454
rect 6840 9302 6960 9330
rect 6840 9194 6868 9302
rect 6987 9276 7295 9285
rect 6987 9274 6993 9276
rect 7049 9274 7073 9276
rect 7129 9274 7153 9276
rect 7209 9274 7233 9276
rect 7289 9274 7295 9276
rect 7049 9222 7051 9274
rect 7231 9222 7233 9274
rect 6987 9220 6993 9222
rect 7049 9220 7073 9222
rect 7129 9220 7153 9222
rect 7209 9220 7233 9222
rect 7289 9220 7295 9222
rect 6987 9211 7295 9220
rect 6840 9166 6960 9194
rect 6932 8838 6960 9166
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 4572 7100 4880 7109
rect 4572 7098 4578 7100
rect 4634 7098 4658 7100
rect 4714 7098 4738 7100
rect 4794 7098 4818 7100
rect 4874 7098 4880 7100
rect 4634 7046 4636 7098
rect 4816 7046 4818 7098
rect 4572 7044 4578 7046
rect 4634 7044 4658 7046
rect 4714 7044 4738 7046
rect 4794 7044 4818 7046
rect 4874 7044 4880 7046
rect 4572 7035 4880 7044
rect 5552 6866 5580 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3344 5778 3372 6190
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5370 4016 5646
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3436 4214 3464 4966
rect 3712 4826 3740 4966
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3738 3372 4082
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3534 3464 4150
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3436 2922 3464 3470
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3712 2854 3740 3470
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3712 2514 3740 2790
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2817 2204 3125 2213
rect 2817 2202 2823 2204
rect 2879 2202 2903 2204
rect 2959 2202 2983 2204
rect 3039 2202 3063 2204
rect 3119 2202 3125 2204
rect 2879 2150 2881 2202
rect 3061 2150 3063 2202
rect 2817 2148 2823 2150
rect 2879 2148 2903 2150
rect 2959 2148 2983 2150
rect 3039 2148 3063 2150
rect 3119 2148 3125 2150
rect 2817 2139 3125 2148
rect 2976 870 3096 898
rect 2976 800 3004 870
rect 2962 0 3018 800
rect 3068 762 3096 870
rect 3252 762 3280 2382
rect 3988 2378 4016 4014
rect 4066 3496 4122 3505
rect 4172 3482 4200 6666
rect 5232 6556 5540 6565
rect 5232 6554 5238 6556
rect 5294 6554 5318 6556
rect 5374 6554 5398 6556
rect 5454 6554 5478 6556
rect 5534 6554 5540 6556
rect 5294 6502 5296 6554
rect 5476 6502 5478 6554
rect 5232 6500 5238 6502
rect 5294 6500 5318 6502
rect 5374 6500 5398 6502
rect 5454 6500 5478 6502
rect 5534 6500 5540 6502
rect 5232 6491 5540 6500
rect 5644 6322 5672 7346
rect 6104 7342 6132 7958
rect 6288 7886 6316 8230
rect 6840 8090 6868 8502
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6987 8188 7295 8197
rect 6987 8186 6993 8188
rect 7049 8186 7073 8188
rect 7129 8186 7153 8188
rect 7209 8186 7233 8188
rect 7289 8186 7295 8188
rect 7049 8134 7051 8186
rect 7231 8134 7233 8186
rect 6987 8132 6993 8134
rect 7049 8132 7073 8134
rect 7129 8132 7153 8134
rect 7209 8132 7233 8134
rect 7289 8132 7295 8134
rect 6987 8123 7295 8132
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6196 6662 6224 7754
rect 6288 7410 6316 7822
rect 6840 7546 6868 8026
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6987 7100 7295 7109
rect 6987 7098 6993 7100
rect 7049 7098 7073 7100
rect 7129 7098 7153 7100
rect 7209 7098 7233 7100
rect 7289 7098 7295 7100
rect 7049 7046 7051 7098
rect 7231 7046 7233 7098
rect 6987 7044 6993 7046
rect 7049 7044 7073 7046
rect 7129 7044 7153 7046
rect 7209 7044 7233 7046
rect 7289 7044 7295 7046
rect 6987 7035 7295 7044
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 4572 6012 4880 6021
rect 4572 6010 4578 6012
rect 4634 6010 4658 6012
rect 4714 6010 4738 6012
rect 4794 6010 4818 6012
rect 4874 6010 4880 6012
rect 4634 5958 4636 6010
rect 4816 5958 4818 6010
rect 4572 5956 4578 5958
rect 4634 5956 4658 5958
rect 4714 5956 4738 5958
rect 4794 5956 4818 5958
rect 4874 5956 4880 5958
rect 4572 5947 4880 5956
rect 4908 5574 4936 6258
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5644 5658 5672 6054
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5644 5630 5764 5658
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 4724 5370 4752 5510
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4572 4924 4880 4933
rect 4572 4922 4578 4924
rect 4634 4922 4658 4924
rect 4714 4922 4738 4924
rect 4794 4922 4818 4924
rect 4874 4922 4880 4924
rect 4634 4870 4636 4922
rect 4816 4870 4818 4922
rect 4572 4868 4578 4870
rect 4634 4868 4658 4870
rect 4714 4868 4738 4870
rect 4794 4868 4818 4870
rect 4874 4868 4880 4870
rect 4572 4859 4880 4868
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4078 4476 4422
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4908 4010 4936 5510
rect 5232 5468 5540 5477
rect 5232 5466 5238 5468
rect 5294 5466 5318 5468
rect 5374 5466 5398 5468
rect 5454 5466 5478 5468
rect 5534 5466 5540 5468
rect 5294 5414 5296 5466
rect 5476 5414 5478 5466
rect 5232 5412 5238 5414
rect 5294 5412 5318 5414
rect 5374 5412 5398 5414
rect 5454 5412 5478 5414
rect 5534 5412 5540 5414
rect 5232 5403 5540 5412
rect 5644 5030 5672 5510
rect 5736 5302 5764 5630
rect 6012 5574 6040 6054
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5370 6040 5510
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5232 4380 5540 4389
rect 5232 4378 5238 4380
rect 5294 4378 5318 4380
rect 5374 4378 5398 4380
rect 5454 4378 5478 4380
rect 5534 4378 5540 4380
rect 5294 4326 5296 4378
rect 5476 4326 5478 4378
rect 5232 4324 5238 4326
rect 5294 4324 5318 4326
rect 5374 4324 5398 4326
rect 5454 4324 5478 4326
rect 5534 4324 5540 4326
rect 5232 4315 5540 4324
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4572 3836 4880 3845
rect 4572 3834 4578 3836
rect 4634 3834 4658 3836
rect 4714 3834 4738 3836
rect 4794 3834 4818 3836
rect 4874 3834 4880 3836
rect 4634 3782 4636 3834
rect 4816 3782 4818 3834
rect 4572 3780 4578 3782
rect 4634 3780 4658 3782
rect 4714 3780 4738 3782
rect 4794 3780 4818 3782
rect 4874 3780 4880 3782
rect 4572 3771 4880 3780
rect 4122 3454 4200 3482
rect 5552 3482 5580 4082
rect 5644 3602 5672 4966
rect 6012 4214 6040 5306
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3738 5764 3878
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5552 3454 5672 3482
rect 6012 3466 6040 4150
rect 4066 3431 4122 3440
rect 5644 3398 5672 3454
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5232 3292 5540 3301
rect 5232 3290 5238 3292
rect 5294 3290 5318 3292
rect 5374 3290 5398 3292
rect 5454 3290 5478 3292
rect 5534 3290 5540 3292
rect 5294 3238 5296 3290
rect 5476 3238 5478 3290
rect 5232 3236 5238 3238
rect 5294 3236 5318 3238
rect 5374 3236 5398 3238
rect 5454 3236 5478 3238
rect 5534 3236 5540 3238
rect 5232 3227 5540 3236
rect 5644 2990 5672 3334
rect 6196 3126 6224 6598
rect 6987 6012 7295 6021
rect 6987 6010 6993 6012
rect 7049 6010 7073 6012
rect 7129 6010 7153 6012
rect 7209 6010 7233 6012
rect 7289 6010 7295 6012
rect 7049 5958 7051 6010
rect 7231 5958 7233 6010
rect 6987 5956 6993 5958
rect 7049 5956 7073 5958
rect 7129 5956 7153 5958
rect 7209 5956 7233 5958
rect 7289 5956 7295 5958
rect 6987 5947 7295 5956
rect 6987 4924 7295 4933
rect 6987 4922 6993 4924
rect 7049 4922 7073 4924
rect 7129 4922 7153 4924
rect 7209 4922 7233 4924
rect 7289 4922 7295 4924
rect 7049 4870 7051 4922
rect 7231 4870 7233 4922
rect 6987 4868 6993 4870
rect 7049 4868 7073 4870
rect 7129 4868 7153 4870
rect 7209 4868 7233 4870
rect 7289 4868 7295 4870
rect 6987 4859 7295 4868
rect 7392 4758 7420 8842
rect 7484 8090 7512 9522
rect 8116 9512 8168 9518
rect 8220 9466 8248 9998
rect 8496 9722 8524 10066
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8168 9460 8248 9466
rect 8116 9454 8248 9460
rect 8128 9438 8248 9454
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7647 8732 7955 8741
rect 7647 8730 7653 8732
rect 7709 8730 7733 8732
rect 7789 8730 7813 8732
rect 7869 8730 7893 8732
rect 7949 8730 7955 8732
rect 7709 8678 7711 8730
rect 7891 8678 7893 8730
rect 7647 8676 7653 8678
rect 7709 8676 7733 8678
rect 7789 8676 7813 8678
rect 7869 8676 7893 8678
rect 7949 8676 7955 8678
rect 7647 8667 7955 8676
rect 8036 8498 8064 8842
rect 8128 8838 8156 9438
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7546 7604 7822
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7647 7644 7955 7653
rect 7647 7642 7653 7644
rect 7709 7642 7733 7644
rect 7789 7642 7813 7644
rect 7869 7642 7893 7644
rect 7949 7642 7955 7644
rect 7709 7590 7711 7642
rect 7891 7590 7893 7642
rect 7647 7588 7653 7590
rect 7709 7588 7733 7590
rect 7789 7588 7813 7590
rect 7869 7588 7893 7590
rect 7949 7588 7955 7590
rect 7647 7579 7955 7588
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6458 7512 6666
rect 7647 6556 7955 6565
rect 7647 6554 7653 6556
rect 7709 6554 7733 6556
rect 7789 6554 7813 6556
rect 7869 6554 7893 6556
rect 7949 6554 7955 6556
rect 7709 6502 7711 6554
rect 7891 6502 7893 6554
rect 7647 6500 7653 6502
rect 7709 6500 7733 6502
rect 7789 6500 7813 6502
rect 7869 6500 7893 6502
rect 7949 6500 7955 6502
rect 7647 6491 7955 6500
rect 8036 6458 8064 7686
rect 8128 7478 8156 8774
rect 8220 8498 8248 9318
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8404 7410 8432 8570
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 7546 8616 7822
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8404 6322 8432 7346
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8496 6118 8524 6598
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7647 5468 7955 5477
rect 7647 5466 7653 5468
rect 7709 5466 7733 5468
rect 7789 5466 7813 5468
rect 7869 5466 7893 5468
rect 7949 5466 7955 5468
rect 7709 5414 7711 5466
rect 7891 5414 7893 5466
rect 7647 5412 7653 5414
rect 7709 5412 7733 5414
rect 7789 5412 7813 5414
rect 7869 5412 7893 5414
rect 7949 5412 7955 5414
rect 7647 5403 7955 5412
rect 8128 4826 8156 5850
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7392 4010 7420 4694
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4146 7512 4558
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 6987 3836 7295 3845
rect 6987 3834 6993 3836
rect 7049 3834 7073 3836
rect 7129 3834 7153 3836
rect 7209 3834 7233 3836
rect 7289 3834 7295 3836
rect 7049 3782 7051 3834
rect 7231 3782 7233 3834
rect 6987 3780 6993 3782
rect 7049 3780 7073 3782
rect 7129 3780 7153 3782
rect 7209 3780 7233 3782
rect 7289 3780 7295 3782
rect 6987 3771 7295 3780
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7300 3126 7328 3334
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 2774 4108 2858
rect 4080 2746 4384 2774
rect 4356 2378 4384 2746
rect 4572 2748 4880 2757
rect 4572 2746 4578 2748
rect 4634 2746 4658 2748
rect 4714 2746 4738 2748
rect 4794 2746 4818 2748
rect 4874 2746 4880 2748
rect 4634 2694 4636 2746
rect 4816 2694 4818 2746
rect 4572 2692 4578 2694
rect 4634 2692 4658 2694
rect 4714 2692 4738 2694
rect 4794 2692 4818 2694
rect 4874 2692 4880 2694
rect 4572 2683 4880 2692
rect 5644 2650 5672 2926
rect 7392 2922 7420 3946
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3738 7512 3878
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 3466 7604 4422
rect 7647 4380 7955 4389
rect 7647 4378 7653 4380
rect 7709 4378 7733 4380
rect 7789 4378 7813 4380
rect 7869 4378 7893 4380
rect 7949 4378 7955 4380
rect 7709 4326 7711 4378
rect 7891 4326 7893 4378
rect 7647 4324 7653 4326
rect 7709 4324 7733 4326
rect 7789 4324 7813 4326
rect 7869 4324 7893 4326
rect 7949 4324 7955 4326
rect 7647 4315 7955 4324
rect 7840 4072 7892 4078
rect 8128 4026 8156 4762
rect 7892 4020 8156 4026
rect 7840 4014 8156 4020
rect 7852 3998 8156 4014
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7760 3738 7788 3878
rect 8220 3754 8248 5510
rect 8496 5166 8524 6054
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 7748 3732 7800 3738
rect 8220 3726 8340 3754
rect 7748 3674 7800 3680
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3058 7512 3334
rect 7647 3292 7955 3301
rect 7647 3290 7653 3292
rect 7709 3290 7733 3292
rect 7789 3290 7813 3292
rect 7869 3290 7893 3292
rect 7949 3290 7955 3292
rect 7709 3238 7711 3290
rect 7891 3238 7893 3290
rect 7647 3236 7653 3238
rect 7709 3236 7733 3238
rect 7789 3236 7813 3238
rect 7869 3236 7893 3238
rect 7949 3236 7955 3238
rect 7647 3227 7955 3236
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 6987 2748 7295 2757
rect 6987 2746 6993 2748
rect 7049 2746 7073 2748
rect 7129 2746 7153 2748
rect 7209 2746 7233 2748
rect 7289 2746 7295 2748
rect 7049 2694 7051 2746
rect 7231 2694 7233 2746
rect 6987 2692 6993 2694
rect 7049 2692 7073 2694
rect 7129 2692 7153 2694
rect 7209 2692 7233 2694
rect 7289 2692 7295 2694
rect 6987 2683 7295 2692
rect 7392 2650 7420 2858
rect 7944 2650 7972 2994
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8220 2446 8248 3606
rect 8312 3194 8340 3726
rect 8496 3602 8524 5102
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8588 4078 8616 4558
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8588 3738 8616 4014
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8312 2582 8340 3130
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 8680 2310 8708 10610
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 9220 10464 9272 10470
rect 10888 10441 10916 10474
rect 9220 10406 9272 10412
rect 10874 10432 10930 10441
rect 9232 10130 9260 10406
rect 9402 10364 9710 10373
rect 10874 10367 10930 10376
rect 9402 10362 9408 10364
rect 9464 10362 9488 10364
rect 9544 10362 9568 10364
rect 9624 10362 9648 10364
rect 9704 10362 9710 10364
rect 9464 10310 9466 10362
rect 9646 10310 9648 10362
rect 9402 10308 9408 10310
rect 9464 10308 9488 10310
rect 9544 10308 9568 10310
rect 9624 10308 9648 10310
rect 9704 10308 9710 10310
rect 9402 10299 9710 10308
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9654 9536 9862
rect 10062 9820 10370 9829
rect 10062 9818 10068 9820
rect 10124 9818 10148 9820
rect 10204 9818 10228 9820
rect 10284 9818 10308 9820
rect 10364 9818 10370 9820
rect 10124 9766 10126 9818
rect 10306 9766 10308 9818
rect 10062 9764 10068 9766
rect 10124 9764 10148 9766
rect 10204 9764 10228 9766
rect 10284 9764 10308 9766
rect 10364 9764 10370 9766
rect 10062 9755 10370 9764
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8634 9076 9454
rect 9402 9276 9710 9285
rect 9402 9274 9408 9276
rect 9464 9274 9488 9276
rect 9544 9274 9568 9276
rect 9624 9274 9648 9276
rect 9704 9274 9710 9276
rect 9464 9222 9466 9274
rect 9646 9222 9648 9274
rect 9402 9220 9408 9222
rect 9464 9220 9488 9222
rect 9544 9220 9568 9222
rect 9624 9220 9648 9222
rect 9704 9220 9710 9222
rect 9402 9211 9710 9220
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7342 9168 7890
rect 9232 7546 9260 8774
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7886 9352 8230
rect 9402 8188 9710 8197
rect 9402 8186 9408 8188
rect 9464 8186 9488 8188
rect 9544 8186 9568 8188
rect 9624 8186 9648 8188
rect 9704 8186 9710 8188
rect 9464 8134 9466 8186
rect 9646 8134 9648 8186
rect 9402 8132 9408 8134
rect 9464 8132 9488 8134
rect 9544 8132 9568 8134
rect 9624 8132 9648 8134
rect 9704 8132 9710 8134
rect 9402 8123 9710 8132
rect 9876 8090 9904 8842
rect 10062 8732 10370 8741
rect 10062 8730 10068 8732
rect 10124 8730 10148 8732
rect 10204 8730 10228 8732
rect 10284 8730 10308 8732
rect 10364 8730 10370 8732
rect 10124 8678 10126 8730
rect 10306 8678 10308 8730
rect 10062 8676 10068 8678
rect 10124 8676 10148 8678
rect 10204 8676 10228 8678
rect 10284 8676 10308 8678
rect 10364 8676 10370 8678
rect 10062 8667 10370 8676
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9402 7100 9710 7109
rect 9402 7098 9408 7100
rect 9464 7098 9488 7100
rect 9544 7098 9568 7100
rect 9624 7098 9648 7100
rect 9704 7098 9710 7100
rect 9464 7046 9466 7098
rect 9646 7046 9648 7098
rect 9402 7044 9408 7046
rect 9464 7044 9488 7046
rect 9544 7044 9568 7046
rect 9624 7044 9648 7046
rect 9704 7044 9710 7046
rect 9402 7035 9710 7044
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9402 6012 9710 6021
rect 9402 6010 9408 6012
rect 9464 6010 9488 6012
rect 9544 6010 9568 6012
rect 9624 6010 9648 6012
rect 9704 6010 9710 6012
rect 9464 5958 9466 6010
rect 9646 5958 9648 6010
rect 9402 5956 9408 5958
rect 9464 5956 9488 5958
rect 9544 5956 9568 5958
rect 9624 5956 9648 5958
rect 9704 5956 9710 5958
rect 9402 5947 9710 5956
rect 9784 5794 9812 7686
rect 9876 7342 9904 7686
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6866 9904 7142
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9968 5914 9996 7686
rect 10062 7644 10370 7653
rect 10062 7642 10068 7644
rect 10124 7642 10148 7644
rect 10204 7642 10228 7644
rect 10284 7642 10308 7644
rect 10364 7642 10370 7644
rect 10124 7590 10126 7642
rect 10306 7590 10308 7642
rect 10062 7588 10068 7590
rect 10124 7588 10148 7590
rect 10204 7588 10228 7590
rect 10284 7588 10308 7590
rect 10364 7588 10370 7590
rect 10062 7579 10370 7588
rect 10428 7410 10456 7686
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10336 6934 10364 7346
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10062 6556 10370 6565
rect 10062 6554 10068 6556
rect 10124 6554 10148 6556
rect 10204 6554 10228 6556
rect 10284 6554 10308 6556
rect 10364 6554 10370 6556
rect 10124 6502 10126 6554
rect 10306 6502 10308 6554
rect 10062 6500 10068 6502
rect 10124 6500 10148 6502
rect 10204 6500 10228 6502
rect 10284 6500 10308 6502
rect 10364 6500 10370 6502
rect 10062 6491 10370 6500
rect 10428 6458 10456 7346
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9784 5766 9904 5794
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4622 8800 4966
rect 8956 4622 8984 5510
rect 9232 5302 9260 5510
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9402 4924 9710 4933
rect 9402 4922 9408 4924
rect 9464 4922 9488 4924
rect 9544 4922 9568 4924
rect 9624 4922 9648 4924
rect 9704 4922 9710 4924
rect 9464 4870 9466 4922
rect 9646 4870 9648 4922
rect 9402 4868 9408 4870
rect 9464 4868 9488 4870
rect 9544 4868 9568 4870
rect 9624 4868 9648 4870
rect 9704 4868 9710 4870
rect 9402 4859 9710 4868
rect 9784 4826 9812 5646
rect 9876 5574 9904 5766
rect 10520 5642 10548 7142
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10062 5468 10370 5477
rect 10062 5466 10068 5468
rect 10124 5466 10148 5468
rect 10204 5466 10228 5468
rect 10284 5466 10308 5468
rect 10364 5466 10370 5468
rect 10124 5414 10126 5466
rect 10306 5414 10308 5466
rect 10062 5412 10068 5414
rect 10124 5412 10148 5414
rect 10204 5412 10228 5414
rect 10284 5412 10308 5414
rect 10364 5412 10370 5414
rect 10062 5403 10370 5412
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4690 9904 4966
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8772 4146 8800 4558
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8772 3534 8800 4082
rect 8956 3942 8984 4558
rect 9876 4146 9904 4626
rect 10062 4380 10370 4389
rect 10062 4378 10068 4380
rect 10124 4378 10148 4380
rect 10204 4378 10228 4380
rect 10284 4378 10308 4380
rect 10364 4378 10370 4380
rect 10124 4326 10126 4378
rect 10306 4326 10308 4378
rect 10062 4324 10068 4326
rect 10124 4324 10148 4326
rect 10204 4324 10228 4326
rect 10284 4324 10308 4326
rect 10364 4324 10370 4326
rect 10062 4315 10370 4324
rect 10612 4146 10640 7890
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9048 3194 9076 4014
rect 9402 3836 9710 3845
rect 9402 3834 9408 3836
rect 9464 3834 9488 3836
rect 9544 3834 9568 3836
rect 9624 3834 9648 3836
rect 9704 3834 9710 3836
rect 9464 3782 9466 3834
rect 9646 3782 9648 3834
rect 9402 3780 9408 3782
rect 9464 3780 9488 3782
rect 9544 3780 9568 3782
rect 9624 3780 9648 3782
rect 9704 3780 9710 3782
rect 9402 3771 9710 3780
rect 9968 3738 9996 4014
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 3194 9904 3402
rect 10062 3292 10370 3301
rect 10062 3290 10068 3292
rect 10124 3290 10148 3292
rect 10204 3290 10228 3292
rect 10284 3290 10308 3292
rect 10364 3290 10370 3292
rect 10124 3238 10126 3290
rect 10306 3238 10308 3290
rect 10062 3236 10068 3238
rect 10124 3236 10148 3238
rect 10204 3236 10228 3238
rect 10284 3236 10308 3238
rect 10364 3236 10370 3238
rect 10062 3227 10370 3236
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9048 2514 9076 3130
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9402 2748 9710 2757
rect 9402 2746 9408 2748
rect 9464 2746 9488 2748
rect 9544 2746 9568 2748
rect 9624 2746 9648 2748
rect 9704 2746 9710 2748
rect 9464 2694 9466 2746
rect 9646 2694 9648 2746
rect 9402 2692 9408 2694
rect 9464 2692 9488 2694
rect 9544 2692 9568 2694
rect 9624 2692 9648 2694
rect 9704 2692 9710 2694
rect 9402 2683 9710 2692
rect 9784 2650 9812 2790
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10428 2514 10456 3674
rect 10704 3194 10732 10202
rect 10874 3360 10930 3369
rect 10874 3295 10930 3304
rect 10888 3194 10916 3295
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 5232 2204 5540 2213
rect 5232 2202 5238 2204
rect 5294 2202 5318 2204
rect 5374 2202 5398 2204
rect 5454 2202 5478 2204
rect 5534 2202 5540 2204
rect 5294 2150 5296 2202
rect 5476 2150 5478 2202
rect 5232 2148 5238 2150
rect 5294 2148 5318 2150
rect 5374 2148 5398 2150
rect 5454 2148 5478 2150
rect 5534 2148 5540 2150
rect 5232 2139 5540 2148
rect 7647 2204 7955 2213
rect 7647 2202 7653 2204
rect 7709 2202 7733 2204
rect 7789 2202 7813 2204
rect 7869 2202 7893 2204
rect 7949 2202 7955 2204
rect 7709 2150 7711 2202
rect 7891 2150 7893 2202
rect 7647 2148 7653 2150
rect 7709 2148 7733 2150
rect 7789 2148 7813 2150
rect 7869 2148 7893 2150
rect 7949 2148 7955 2150
rect 7647 2139 7955 2148
rect 8772 1306 8800 2314
rect 10062 2204 10370 2213
rect 10062 2202 10068 2204
rect 10124 2202 10148 2204
rect 10204 2202 10228 2204
rect 10284 2202 10308 2204
rect 10364 2202 10370 2204
rect 10124 2150 10126 2202
rect 10306 2150 10308 2202
rect 10062 2148 10068 2150
rect 10124 2148 10148 2150
rect 10204 2148 10228 2150
rect 10284 2148 10308 2150
rect 10364 2148 10370 2150
rect 10062 2139 10370 2148
rect 8772 1278 8984 1306
rect 8956 800 8984 1278
rect 3068 734 3280 762
rect 8942 0 8998 800
<< via2 >>
rect 2163 11450 2219 11452
rect 2243 11450 2299 11452
rect 2323 11450 2379 11452
rect 2403 11450 2459 11452
rect 2163 11398 2209 11450
rect 2209 11398 2219 11450
rect 2243 11398 2273 11450
rect 2273 11398 2285 11450
rect 2285 11398 2299 11450
rect 2323 11398 2337 11450
rect 2337 11398 2349 11450
rect 2349 11398 2379 11450
rect 2403 11398 2413 11450
rect 2413 11398 2459 11450
rect 2163 11396 2219 11398
rect 2243 11396 2299 11398
rect 2323 11396 2379 11398
rect 2403 11396 2459 11398
rect 4578 11450 4634 11452
rect 4658 11450 4714 11452
rect 4738 11450 4794 11452
rect 4818 11450 4874 11452
rect 4578 11398 4624 11450
rect 4624 11398 4634 11450
rect 4658 11398 4688 11450
rect 4688 11398 4700 11450
rect 4700 11398 4714 11450
rect 4738 11398 4752 11450
rect 4752 11398 4764 11450
rect 4764 11398 4794 11450
rect 4818 11398 4828 11450
rect 4828 11398 4874 11450
rect 4578 11396 4634 11398
rect 4658 11396 4714 11398
rect 4738 11396 4794 11398
rect 4818 11396 4874 11398
rect 6993 11450 7049 11452
rect 7073 11450 7129 11452
rect 7153 11450 7209 11452
rect 7233 11450 7289 11452
rect 6993 11398 7039 11450
rect 7039 11398 7049 11450
rect 7073 11398 7103 11450
rect 7103 11398 7115 11450
rect 7115 11398 7129 11450
rect 7153 11398 7167 11450
rect 7167 11398 7179 11450
rect 7179 11398 7209 11450
rect 7233 11398 7243 11450
rect 7243 11398 7289 11450
rect 6993 11396 7049 11398
rect 7073 11396 7129 11398
rect 7153 11396 7209 11398
rect 7233 11396 7289 11398
rect 9408 11450 9464 11452
rect 9488 11450 9544 11452
rect 9568 11450 9624 11452
rect 9648 11450 9704 11452
rect 9408 11398 9454 11450
rect 9454 11398 9464 11450
rect 9488 11398 9518 11450
rect 9518 11398 9530 11450
rect 9530 11398 9544 11450
rect 9568 11398 9582 11450
rect 9582 11398 9594 11450
rect 9594 11398 9624 11450
rect 9648 11398 9658 11450
rect 9658 11398 9704 11450
rect 9408 11396 9464 11398
rect 9488 11396 9544 11398
rect 9568 11396 9624 11398
rect 9648 11396 9704 11398
rect 2823 10906 2879 10908
rect 2903 10906 2959 10908
rect 2983 10906 3039 10908
rect 3063 10906 3119 10908
rect 2823 10854 2869 10906
rect 2869 10854 2879 10906
rect 2903 10854 2933 10906
rect 2933 10854 2945 10906
rect 2945 10854 2959 10906
rect 2983 10854 2997 10906
rect 2997 10854 3009 10906
rect 3009 10854 3039 10906
rect 3063 10854 3073 10906
rect 3073 10854 3119 10906
rect 2823 10852 2879 10854
rect 2903 10852 2959 10854
rect 2983 10852 3039 10854
rect 3063 10852 3119 10854
rect 938 10376 994 10432
rect 2163 10362 2219 10364
rect 2243 10362 2299 10364
rect 2323 10362 2379 10364
rect 2403 10362 2459 10364
rect 2163 10310 2209 10362
rect 2209 10310 2219 10362
rect 2243 10310 2273 10362
rect 2273 10310 2285 10362
rect 2285 10310 2299 10362
rect 2323 10310 2337 10362
rect 2337 10310 2349 10362
rect 2349 10310 2379 10362
rect 2403 10310 2413 10362
rect 2413 10310 2459 10362
rect 2163 10308 2219 10310
rect 2243 10308 2299 10310
rect 2323 10308 2379 10310
rect 2403 10308 2459 10310
rect 5238 10906 5294 10908
rect 5318 10906 5374 10908
rect 5398 10906 5454 10908
rect 5478 10906 5534 10908
rect 5238 10854 5284 10906
rect 5284 10854 5294 10906
rect 5318 10854 5348 10906
rect 5348 10854 5360 10906
rect 5360 10854 5374 10906
rect 5398 10854 5412 10906
rect 5412 10854 5424 10906
rect 5424 10854 5454 10906
rect 5478 10854 5488 10906
rect 5488 10854 5534 10906
rect 5238 10852 5294 10854
rect 5318 10852 5374 10854
rect 5398 10852 5454 10854
rect 5478 10852 5534 10854
rect 2823 9818 2879 9820
rect 2903 9818 2959 9820
rect 2983 9818 3039 9820
rect 3063 9818 3119 9820
rect 2823 9766 2869 9818
rect 2869 9766 2879 9818
rect 2903 9766 2933 9818
rect 2933 9766 2945 9818
rect 2945 9766 2959 9818
rect 2983 9766 2997 9818
rect 2997 9766 3009 9818
rect 3009 9766 3039 9818
rect 3063 9766 3073 9818
rect 3073 9766 3119 9818
rect 2823 9764 2879 9766
rect 2903 9764 2959 9766
rect 2983 9764 3039 9766
rect 3063 9764 3119 9766
rect 2163 9274 2219 9276
rect 2243 9274 2299 9276
rect 2323 9274 2379 9276
rect 2403 9274 2459 9276
rect 2163 9222 2209 9274
rect 2209 9222 2219 9274
rect 2243 9222 2273 9274
rect 2273 9222 2285 9274
rect 2285 9222 2299 9274
rect 2323 9222 2337 9274
rect 2337 9222 2349 9274
rect 2349 9222 2379 9274
rect 2403 9222 2413 9274
rect 2413 9222 2459 9274
rect 2163 9220 2219 9222
rect 2243 9220 2299 9222
rect 2323 9220 2379 9222
rect 2403 9220 2459 9222
rect 2163 8186 2219 8188
rect 2243 8186 2299 8188
rect 2323 8186 2379 8188
rect 2403 8186 2459 8188
rect 2163 8134 2209 8186
rect 2209 8134 2219 8186
rect 2243 8134 2273 8186
rect 2273 8134 2285 8186
rect 2285 8134 2299 8186
rect 2323 8134 2337 8186
rect 2337 8134 2349 8186
rect 2349 8134 2379 8186
rect 2403 8134 2413 8186
rect 2413 8134 2459 8186
rect 2163 8132 2219 8134
rect 2243 8132 2299 8134
rect 2323 8132 2379 8134
rect 2403 8132 2459 8134
rect 2823 8730 2879 8732
rect 2903 8730 2959 8732
rect 2983 8730 3039 8732
rect 3063 8730 3119 8732
rect 2823 8678 2869 8730
rect 2869 8678 2879 8730
rect 2903 8678 2933 8730
rect 2933 8678 2945 8730
rect 2945 8678 2959 8730
rect 2983 8678 2997 8730
rect 2997 8678 3009 8730
rect 3009 8678 3039 8730
rect 3063 8678 3073 8730
rect 3073 8678 3119 8730
rect 2823 8676 2879 8678
rect 2903 8676 2959 8678
rect 2983 8676 3039 8678
rect 3063 8676 3119 8678
rect 2823 7642 2879 7644
rect 2903 7642 2959 7644
rect 2983 7642 3039 7644
rect 3063 7642 3119 7644
rect 2823 7590 2869 7642
rect 2869 7590 2879 7642
rect 2903 7590 2933 7642
rect 2933 7590 2945 7642
rect 2945 7590 2959 7642
rect 2983 7590 2997 7642
rect 2997 7590 3009 7642
rect 3009 7590 3039 7642
rect 3063 7590 3073 7642
rect 3073 7590 3119 7642
rect 2823 7588 2879 7590
rect 2903 7588 2959 7590
rect 2983 7588 3039 7590
rect 3063 7588 3119 7590
rect 2163 7098 2219 7100
rect 2243 7098 2299 7100
rect 2323 7098 2379 7100
rect 2403 7098 2459 7100
rect 2163 7046 2209 7098
rect 2209 7046 2219 7098
rect 2243 7046 2273 7098
rect 2273 7046 2285 7098
rect 2285 7046 2299 7098
rect 2323 7046 2337 7098
rect 2337 7046 2349 7098
rect 2349 7046 2379 7098
rect 2403 7046 2413 7098
rect 2413 7046 2459 7098
rect 2163 7044 2219 7046
rect 2243 7044 2299 7046
rect 2323 7044 2379 7046
rect 2403 7044 2459 7046
rect 2823 6554 2879 6556
rect 2903 6554 2959 6556
rect 2983 6554 3039 6556
rect 3063 6554 3119 6556
rect 2823 6502 2869 6554
rect 2869 6502 2879 6554
rect 2903 6502 2933 6554
rect 2933 6502 2945 6554
rect 2945 6502 2959 6554
rect 2983 6502 2997 6554
rect 2997 6502 3009 6554
rect 3009 6502 3039 6554
rect 3063 6502 3073 6554
rect 3073 6502 3119 6554
rect 2823 6500 2879 6502
rect 2903 6500 2959 6502
rect 2983 6500 3039 6502
rect 3063 6500 3119 6502
rect 2163 6010 2219 6012
rect 2243 6010 2299 6012
rect 2323 6010 2379 6012
rect 2403 6010 2459 6012
rect 2163 5958 2209 6010
rect 2209 5958 2219 6010
rect 2243 5958 2273 6010
rect 2273 5958 2285 6010
rect 2285 5958 2299 6010
rect 2323 5958 2337 6010
rect 2337 5958 2349 6010
rect 2349 5958 2379 6010
rect 2403 5958 2413 6010
rect 2413 5958 2459 6010
rect 2163 5956 2219 5958
rect 2243 5956 2299 5958
rect 2323 5956 2379 5958
rect 2403 5956 2459 5958
rect 2823 5466 2879 5468
rect 2903 5466 2959 5468
rect 2983 5466 3039 5468
rect 3063 5466 3119 5468
rect 2823 5414 2869 5466
rect 2869 5414 2879 5466
rect 2903 5414 2933 5466
rect 2933 5414 2945 5466
rect 2945 5414 2959 5466
rect 2983 5414 2997 5466
rect 2997 5414 3009 5466
rect 3009 5414 3039 5466
rect 3063 5414 3073 5466
rect 3073 5414 3119 5466
rect 2823 5412 2879 5414
rect 2903 5412 2959 5414
rect 2983 5412 3039 5414
rect 3063 5412 3119 5414
rect 2163 4922 2219 4924
rect 2243 4922 2299 4924
rect 2323 4922 2379 4924
rect 2403 4922 2459 4924
rect 2163 4870 2209 4922
rect 2209 4870 2219 4922
rect 2243 4870 2273 4922
rect 2273 4870 2285 4922
rect 2285 4870 2299 4922
rect 2323 4870 2337 4922
rect 2337 4870 2349 4922
rect 2349 4870 2379 4922
rect 2403 4870 2413 4922
rect 2413 4870 2459 4922
rect 2163 4868 2219 4870
rect 2243 4868 2299 4870
rect 2323 4868 2379 4870
rect 2403 4868 2459 4870
rect 2823 4378 2879 4380
rect 2903 4378 2959 4380
rect 2983 4378 3039 4380
rect 3063 4378 3119 4380
rect 2823 4326 2869 4378
rect 2869 4326 2879 4378
rect 2903 4326 2933 4378
rect 2933 4326 2945 4378
rect 2945 4326 2959 4378
rect 2983 4326 2997 4378
rect 2997 4326 3009 4378
rect 3009 4326 3039 4378
rect 3063 4326 3073 4378
rect 3073 4326 3119 4378
rect 2823 4324 2879 4326
rect 2903 4324 2959 4326
rect 2983 4324 3039 4326
rect 3063 4324 3119 4326
rect 2163 3834 2219 3836
rect 2243 3834 2299 3836
rect 2323 3834 2379 3836
rect 2403 3834 2459 3836
rect 2163 3782 2209 3834
rect 2209 3782 2219 3834
rect 2243 3782 2273 3834
rect 2273 3782 2285 3834
rect 2285 3782 2299 3834
rect 2323 3782 2337 3834
rect 2337 3782 2349 3834
rect 2349 3782 2379 3834
rect 2403 3782 2413 3834
rect 2413 3782 2459 3834
rect 2163 3780 2219 3782
rect 2243 3780 2299 3782
rect 2323 3780 2379 3782
rect 2403 3780 2459 3782
rect 2823 3290 2879 3292
rect 2903 3290 2959 3292
rect 2983 3290 3039 3292
rect 3063 3290 3119 3292
rect 2823 3238 2869 3290
rect 2869 3238 2879 3290
rect 2903 3238 2933 3290
rect 2933 3238 2945 3290
rect 2945 3238 2959 3290
rect 2983 3238 2997 3290
rect 2997 3238 3009 3290
rect 3009 3238 3039 3290
rect 3063 3238 3073 3290
rect 3073 3238 3119 3290
rect 2823 3236 2879 3238
rect 2903 3236 2959 3238
rect 2983 3236 3039 3238
rect 3063 3236 3119 3238
rect 2163 2746 2219 2748
rect 2243 2746 2299 2748
rect 2323 2746 2379 2748
rect 2403 2746 2459 2748
rect 2163 2694 2209 2746
rect 2209 2694 2219 2746
rect 2243 2694 2273 2746
rect 2273 2694 2285 2746
rect 2285 2694 2299 2746
rect 2323 2694 2337 2746
rect 2337 2694 2349 2746
rect 2349 2694 2379 2746
rect 2403 2694 2413 2746
rect 2413 2694 2459 2746
rect 2163 2692 2219 2694
rect 2243 2692 2299 2694
rect 2323 2692 2379 2694
rect 2403 2692 2459 2694
rect 4578 10362 4634 10364
rect 4658 10362 4714 10364
rect 4738 10362 4794 10364
rect 4818 10362 4874 10364
rect 4578 10310 4624 10362
rect 4624 10310 4634 10362
rect 4658 10310 4688 10362
rect 4688 10310 4700 10362
rect 4700 10310 4714 10362
rect 4738 10310 4752 10362
rect 4752 10310 4764 10362
rect 4764 10310 4794 10362
rect 4818 10310 4828 10362
rect 4828 10310 4874 10362
rect 4578 10308 4634 10310
rect 4658 10308 4714 10310
rect 4738 10308 4794 10310
rect 4818 10308 4874 10310
rect 5238 9818 5294 9820
rect 5318 9818 5374 9820
rect 5398 9818 5454 9820
rect 5478 9818 5534 9820
rect 5238 9766 5284 9818
rect 5284 9766 5294 9818
rect 5318 9766 5348 9818
rect 5348 9766 5360 9818
rect 5360 9766 5374 9818
rect 5398 9766 5412 9818
rect 5412 9766 5424 9818
rect 5424 9766 5454 9818
rect 5478 9766 5488 9818
rect 5488 9766 5534 9818
rect 5238 9764 5294 9766
rect 5318 9764 5374 9766
rect 5398 9764 5454 9766
rect 5478 9764 5534 9766
rect 6993 10362 7049 10364
rect 7073 10362 7129 10364
rect 7153 10362 7209 10364
rect 7233 10362 7289 10364
rect 6993 10310 7039 10362
rect 7039 10310 7049 10362
rect 7073 10310 7103 10362
rect 7103 10310 7115 10362
rect 7115 10310 7129 10362
rect 7153 10310 7167 10362
rect 7167 10310 7179 10362
rect 7179 10310 7209 10362
rect 7233 10310 7243 10362
rect 7243 10310 7289 10362
rect 6993 10308 7049 10310
rect 7073 10308 7129 10310
rect 7153 10308 7209 10310
rect 7233 10308 7289 10310
rect 4578 9274 4634 9276
rect 4658 9274 4714 9276
rect 4738 9274 4794 9276
rect 4818 9274 4874 9276
rect 4578 9222 4624 9274
rect 4624 9222 4634 9274
rect 4658 9222 4688 9274
rect 4688 9222 4700 9274
rect 4700 9222 4714 9274
rect 4738 9222 4752 9274
rect 4752 9222 4764 9274
rect 4764 9222 4794 9274
rect 4818 9222 4828 9274
rect 4828 9222 4874 9274
rect 4578 9220 4634 9222
rect 4658 9220 4714 9222
rect 4738 9220 4794 9222
rect 4818 9220 4874 9222
rect 5238 8730 5294 8732
rect 5318 8730 5374 8732
rect 5398 8730 5454 8732
rect 5478 8730 5534 8732
rect 5238 8678 5284 8730
rect 5284 8678 5294 8730
rect 5318 8678 5348 8730
rect 5348 8678 5360 8730
rect 5360 8678 5374 8730
rect 5398 8678 5412 8730
rect 5412 8678 5424 8730
rect 5424 8678 5454 8730
rect 5478 8678 5488 8730
rect 5488 8678 5534 8730
rect 5238 8676 5294 8678
rect 5318 8676 5374 8678
rect 5398 8676 5454 8678
rect 5478 8676 5534 8678
rect 4578 8186 4634 8188
rect 4658 8186 4714 8188
rect 4738 8186 4794 8188
rect 4818 8186 4874 8188
rect 4578 8134 4624 8186
rect 4624 8134 4634 8186
rect 4658 8134 4688 8186
rect 4688 8134 4700 8186
rect 4700 8134 4714 8186
rect 4738 8134 4752 8186
rect 4752 8134 4764 8186
rect 4764 8134 4794 8186
rect 4818 8134 4828 8186
rect 4828 8134 4874 8186
rect 4578 8132 4634 8134
rect 4658 8132 4714 8134
rect 4738 8132 4794 8134
rect 4818 8132 4874 8134
rect 5238 7642 5294 7644
rect 5318 7642 5374 7644
rect 5398 7642 5454 7644
rect 5478 7642 5534 7644
rect 5238 7590 5284 7642
rect 5284 7590 5294 7642
rect 5318 7590 5348 7642
rect 5348 7590 5360 7642
rect 5360 7590 5374 7642
rect 5398 7590 5412 7642
rect 5412 7590 5424 7642
rect 5424 7590 5454 7642
rect 5478 7590 5488 7642
rect 5488 7590 5534 7642
rect 5238 7588 5294 7590
rect 5318 7588 5374 7590
rect 5398 7588 5454 7590
rect 5478 7588 5534 7590
rect 7653 10906 7709 10908
rect 7733 10906 7789 10908
rect 7813 10906 7869 10908
rect 7893 10906 7949 10908
rect 7653 10854 7699 10906
rect 7699 10854 7709 10906
rect 7733 10854 7763 10906
rect 7763 10854 7775 10906
rect 7775 10854 7789 10906
rect 7813 10854 7827 10906
rect 7827 10854 7839 10906
rect 7839 10854 7869 10906
rect 7893 10854 7903 10906
rect 7903 10854 7949 10906
rect 7653 10852 7709 10854
rect 7733 10852 7789 10854
rect 7813 10852 7869 10854
rect 7893 10852 7949 10854
rect 7653 9818 7709 9820
rect 7733 9818 7789 9820
rect 7813 9818 7869 9820
rect 7893 9818 7949 9820
rect 7653 9766 7699 9818
rect 7699 9766 7709 9818
rect 7733 9766 7763 9818
rect 7763 9766 7775 9818
rect 7775 9766 7789 9818
rect 7813 9766 7827 9818
rect 7827 9766 7839 9818
rect 7839 9766 7869 9818
rect 7893 9766 7903 9818
rect 7903 9766 7949 9818
rect 7653 9764 7709 9766
rect 7733 9764 7789 9766
rect 7813 9764 7869 9766
rect 7893 9764 7949 9766
rect 10068 10906 10124 10908
rect 10148 10906 10204 10908
rect 10228 10906 10284 10908
rect 10308 10906 10364 10908
rect 10068 10854 10114 10906
rect 10114 10854 10124 10906
rect 10148 10854 10178 10906
rect 10178 10854 10190 10906
rect 10190 10854 10204 10906
rect 10228 10854 10242 10906
rect 10242 10854 10254 10906
rect 10254 10854 10284 10906
rect 10308 10854 10318 10906
rect 10318 10854 10364 10906
rect 10068 10852 10124 10854
rect 10148 10852 10204 10854
rect 10228 10852 10284 10854
rect 10308 10852 10364 10854
rect 6993 9274 7049 9276
rect 7073 9274 7129 9276
rect 7153 9274 7209 9276
rect 7233 9274 7289 9276
rect 6993 9222 7039 9274
rect 7039 9222 7049 9274
rect 7073 9222 7103 9274
rect 7103 9222 7115 9274
rect 7115 9222 7129 9274
rect 7153 9222 7167 9274
rect 7167 9222 7179 9274
rect 7179 9222 7209 9274
rect 7233 9222 7243 9274
rect 7243 9222 7289 9274
rect 6993 9220 7049 9222
rect 7073 9220 7129 9222
rect 7153 9220 7209 9222
rect 7233 9220 7289 9222
rect 4578 7098 4634 7100
rect 4658 7098 4714 7100
rect 4738 7098 4794 7100
rect 4818 7098 4874 7100
rect 4578 7046 4624 7098
rect 4624 7046 4634 7098
rect 4658 7046 4688 7098
rect 4688 7046 4700 7098
rect 4700 7046 4714 7098
rect 4738 7046 4752 7098
rect 4752 7046 4764 7098
rect 4764 7046 4794 7098
rect 4818 7046 4828 7098
rect 4828 7046 4874 7098
rect 4578 7044 4634 7046
rect 4658 7044 4714 7046
rect 4738 7044 4794 7046
rect 4818 7044 4874 7046
rect 2823 2202 2879 2204
rect 2903 2202 2959 2204
rect 2983 2202 3039 2204
rect 3063 2202 3119 2204
rect 2823 2150 2869 2202
rect 2869 2150 2879 2202
rect 2903 2150 2933 2202
rect 2933 2150 2945 2202
rect 2945 2150 2959 2202
rect 2983 2150 2997 2202
rect 2997 2150 3009 2202
rect 3009 2150 3039 2202
rect 3063 2150 3073 2202
rect 3073 2150 3119 2202
rect 2823 2148 2879 2150
rect 2903 2148 2959 2150
rect 2983 2148 3039 2150
rect 3063 2148 3119 2150
rect 4066 3440 4122 3496
rect 5238 6554 5294 6556
rect 5318 6554 5374 6556
rect 5398 6554 5454 6556
rect 5478 6554 5534 6556
rect 5238 6502 5284 6554
rect 5284 6502 5294 6554
rect 5318 6502 5348 6554
rect 5348 6502 5360 6554
rect 5360 6502 5374 6554
rect 5398 6502 5412 6554
rect 5412 6502 5424 6554
rect 5424 6502 5454 6554
rect 5478 6502 5488 6554
rect 5488 6502 5534 6554
rect 5238 6500 5294 6502
rect 5318 6500 5374 6502
rect 5398 6500 5454 6502
rect 5478 6500 5534 6502
rect 6993 8186 7049 8188
rect 7073 8186 7129 8188
rect 7153 8186 7209 8188
rect 7233 8186 7289 8188
rect 6993 8134 7039 8186
rect 7039 8134 7049 8186
rect 7073 8134 7103 8186
rect 7103 8134 7115 8186
rect 7115 8134 7129 8186
rect 7153 8134 7167 8186
rect 7167 8134 7179 8186
rect 7179 8134 7209 8186
rect 7233 8134 7243 8186
rect 7243 8134 7289 8186
rect 6993 8132 7049 8134
rect 7073 8132 7129 8134
rect 7153 8132 7209 8134
rect 7233 8132 7289 8134
rect 6993 7098 7049 7100
rect 7073 7098 7129 7100
rect 7153 7098 7209 7100
rect 7233 7098 7289 7100
rect 6993 7046 7039 7098
rect 7039 7046 7049 7098
rect 7073 7046 7103 7098
rect 7103 7046 7115 7098
rect 7115 7046 7129 7098
rect 7153 7046 7167 7098
rect 7167 7046 7179 7098
rect 7179 7046 7209 7098
rect 7233 7046 7243 7098
rect 7243 7046 7289 7098
rect 6993 7044 7049 7046
rect 7073 7044 7129 7046
rect 7153 7044 7209 7046
rect 7233 7044 7289 7046
rect 4578 6010 4634 6012
rect 4658 6010 4714 6012
rect 4738 6010 4794 6012
rect 4818 6010 4874 6012
rect 4578 5958 4624 6010
rect 4624 5958 4634 6010
rect 4658 5958 4688 6010
rect 4688 5958 4700 6010
rect 4700 5958 4714 6010
rect 4738 5958 4752 6010
rect 4752 5958 4764 6010
rect 4764 5958 4794 6010
rect 4818 5958 4828 6010
rect 4828 5958 4874 6010
rect 4578 5956 4634 5958
rect 4658 5956 4714 5958
rect 4738 5956 4794 5958
rect 4818 5956 4874 5958
rect 4578 4922 4634 4924
rect 4658 4922 4714 4924
rect 4738 4922 4794 4924
rect 4818 4922 4874 4924
rect 4578 4870 4624 4922
rect 4624 4870 4634 4922
rect 4658 4870 4688 4922
rect 4688 4870 4700 4922
rect 4700 4870 4714 4922
rect 4738 4870 4752 4922
rect 4752 4870 4764 4922
rect 4764 4870 4794 4922
rect 4818 4870 4828 4922
rect 4828 4870 4874 4922
rect 4578 4868 4634 4870
rect 4658 4868 4714 4870
rect 4738 4868 4794 4870
rect 4818 4868 4874 4870
rect 5238 5466 5294 5468
rect 5318 5466 5374 5468
rect 5398 5466 5454 5468
rect 5478 5466 5534 5468
rect 5238 5414 5284 5466
rect 5284 5414 5294 5466
rect 5318 5414 5348 5466
rect 5348 5414 5360 5466
rect 5360 5414 5374 5466
rect 5398 5414 5412 5466
rect 5412 5414 5424 5466
rect 5424 5414 5454 5466
rect 5478 5414 5488 5466
rect 5488 5414 5534 5466
rect 5238 5412 5294 5414
rect 5318 5412 5374 5414
rect 5398 5412 5454 5414
rect 5478 5412 5534 5414
rect 5238 4378 5294 4380
rect 5318 4378 5374 4380
rect 5398 4378 5454 4380
rect 5478 4378 5534 4380
rect 5238 4326 5284 4378
rect 5284 4326 5294 4378
rect 5318 4326 5348 4378
rect 5348 4326 5360 4378
rect 5360 4326 5374 4378
rect 5398 4326 5412 4378
rect 5412 4326 5424 4378
rect 5424 4326 5454 4378
rect 5478 4326 5488 4378
rect 5488 4326 5534 4378
rect 5238 4324 5294 4326
rect 5318 4324 5374 4326
rect 5398 4324 5454 4326
rect 5478 4324 5534 4326
rect 4578 3834 4634 3836
rect 4658 3834 4714 3836
rect 4738 3834 4794 3836
rect 4818 3834 4874 3836
rect 4578 3782 4624 3834
rect 4624 3782 4634 3834
rect 4658 3782 4688 3834
rect 4688 3782 4700 3834
rect 4700 3782 4714 3834
rect 4738 3782 4752 3834
rect 4752 3782 4764 3834
rect 4764 3782 4794 3834
rect 4818 3782 4828 3834
rect 4828 3782 4874 3834
rect 4578 3780 4634 3782
rect 4658 3780 4714 3782
rect 4738 3780 4794 3782
rect 4818 3780 4874 3782
rect 5238 3290 5294 3292
rect 5318 3290 5374 3292
rect 5398 3290 5454 3292
rect 5478 3290 5534 3292
rect 5238 3238 5284 3290
rect 5284 3238 5294 3290
rect 5318 3238 5348 3290
rect 5348 3238 5360 3290
rect 5360 3238 5374 3290
rect 5398 3238 5412 3290
rect 5412 3238 5424 3290
rect 5424 3238 5454 3290
rect 5478 3238 5488 3290
rect 5488 3238 5534 3290
rect 5238 3236 5294 3238
rect 5318 3236 5374 3238
rect 5398 3236 5454 3238
rect 5478 3236 5534 3238
rect 6993 6010 7049 6012
rect 7073 6010 7129 6012
rect 7153 6010 7209 6012
rect 7233 6010 7289 6012
rect 6993 5958 7039 6010
rect 7039 5958 7049 6010
rect 7073 5958 7103 6010
rect 7103 5958 7115 6010
rect 7115 5958 7129 6010
rect 7153 5958 7167 6010
rect 7167 5958 7179 6010
rect 7179 5958 7209 6010
rect 7233 5958 7243 6010
rect 7243 5958 7289 6010
rect 6993 5956 7049 5958
rect 7073 5956 7129 5958
rect 7153 5956 7209 5958
rect 7233 5956 7289 5958
rect 6993 4922 7049 4924
rect 7073 4922 7129 4924
rect 7153 4922 7209 4924
rect 7233 4922 7289 4924
rect 6993 4870 7039 4922
rect 7039 4870 7049 4922
rect 7073 4870 7103 4922
rect 7103 4870 7115 4922
rect 7115 4870 7129 4922
rect 7153 4870 7167 4922
rect 7167 4870 7179 4922
rect 7179 4870 7209 4922
rect 7233 4870 7243 4922
rect 7243 4870 7289 4922
rect 6993 4868 7049 4870
rect 7073 4868 7129 4870
rect 7153 4868 7209 4870
rect 7233 4868 7289 4870
rect 7653 8730 7709 8732
rect 7733 8730 7789 8732
rect 7813 8730 7869 8732
rect 7893 8730 7949 8732
rect 7653 8678 7699 8730
rect 7699 8678 7709 8730
rect 7733 8678 7763 8730
rect 7763 8678 7775 8730
rect 7775 8678 7789 8730
rect 7813 8678 7827 8730
rect 7827 8678 7839 8730
rect 7839 8678 7869 8730
rect 7893 8678 7903 8730
rect 7903 8678 7949 8730
rect 7653 8676 7709 8678
rect 7733 8676 7789 8678
rect 7813 8676 7869 8678
rect 7893 8676 7949 8678
rect 7653 7642 7709 7644
rect 7733 7642 7789 7644
rect 7813 7642 7869 7644
rect 7893 7642 7949 7644
rect 7653 7590 7699 7642
rect 7699 7590 7709 7642
rect 7733 7590 7763 7642
rect 7763 7590 7775 7642
rect 7775 7590 7789 7642
rect 7813 7590 7827 7642
rect 7827 7590 7839 7642
rect 7839 7590 7869 7642
rect 7893 7590 7903 7642
rect 7903 7590 7949 7642
rect 7653 7588 7709 7590
rect 7733 7588 7789 7590
rect 7813 7588 7869 7590
rect 7893 7588 7949 7590
rect 7653 6554 7709 6556
rect 7733 6554 7789 6556
rect 7813 6554 7869 6556
rect 7893 6554 7949 6556
rect 7653 6502 7699 6554
rect 7699 6502 7709 6554
rect 7733 6502 7763 6554
rect 7763 6502 7775 6554
rect 7775 6502 7789 6554
rect 7813 6502 7827 6554
rect 7827 6502 7839 6554
rect 7839 6502 7869 6554
rect 7893 6502 7903 6554
rect 7903 6502 7949 6554
rect 7653 6500 7709 6502
rect 7733 6500 7789 6502
rect 7813 6500 7869 6502
rect 7893 6500 7949 6502
rect 7653 5466 7709 5468
rect 7733 5466 7789 5468
rect 7813 5466 7869 5468
rect 7893 5466 7949 5468
rect 7653 5414 7699 5466
rect 7699 5414 7709 5466
rect 7733 5414 7763 5466
rect 7763 5414 7775 5466
rect 7775 5414 7789 5466
rect 7813 5414 7827 5466
rect 7827 5414 7839 5466
rect 7839 5414 7869 5466
rect 7893 5414 7903 5466
rect 7903 5414 7949 5466
rect 7653 5412 7709 5414
rect 7733 5412 7789 5414
rect 7813 5412 7869 5414
rect 7893 5412 7949 5414
rect 6993 3834 7049 3836
rect 7073 3834 7129 3836
rect 7153 3834 7209 3836
rect 7233 3834 7289 3836
rect 6993 3782 7039 3834
rect 7039 3782 7049 3834
rect 7073 3782 7103 3834
rect 7103 3782 7115 3834
rect 7115 3782 7129 3834
rect 7153 3782 7167 3834
rect 7167 3782 7179 3834
rect 7179 3782 7209 3834
rect 7233 3782 7243 3834
rect 7243 3782 7289 3834
rect 6993 3780 7049 3782
rect 7073 3780 7129 3782
rect 7153 3780 7209 3782
rect 7233 3780 7289 3782
rect 4578 2746 4634 2748
rect 4658 2746 4714 2748
rect 4738 2746 4794 2748
rect 4818 2746 4874 2748
rect 4578 2694 4624 2746
rect 4624 2694 4634 2746
rect 4658 2694 4688 2746
rect 4688 2694 4700 2746
rect 4700 2694 4714 2746
rect 4738 2694 4752 2746
rect 4752 2694 4764 2746
rect 4764 2694 4794 2746
rect 4818 2694 4828 2746
rect 4828 2694 4874 2746
rect 4578 2692 4634 2694
rect 4658 2692 4714 2694
rect 4738 2692 4794 2694
rect 4818 2692 4874 2694
rect 7653 4378 7709 4380
rect 7733 4378 7789 4380
rect 7813 4378 7869 4380
rect 7893 4378 7949 4380
rect 7653 4326 7699 4378
rect 7699 4326 7709 4378
rect 7733 4326 7763 4378
rect 7763 4326 7775 4378
rect 7775 4326 7789 4378
rect 7813 4326 7827 4378
rect 7827 4326 7839 4378
rect 7839 4326 7869 4378
rect 7893 4326 7903 4378
rect 7903 4326 7949 4378
rect 7653 4324 7709 4326
rect 7733 4324 7789 4326
rect 7813 4324 7869 4326
rect 7893 4324 7949 4326
rect 7653 3290 7709 3292
rect 7733 3290 7789 3292
rect 7813 3290 7869 3292
rect 7893 3290 7949 3292
rect 7653 3238 7699 3290
rect 7699 3238 7709 3290
rect 7733 3238 7763 3290
rect 7763 3238 7775 3290
rect 7775 3238 7789 3290
rect 7813 3238 7827 3290
rect 7827 3238 7839 3290
rect 7839 3238 7869 3290
rect 7893 3238 7903 3290
rect 7903 3238 7949 3290
rect 7653 3236 7709 3238
rect 7733 3236 7789 3238
rect 7813 3236 7869 3238
rect 7893 3236 7949 3238
rect 6993 2746 7049 2748
rect 7073 2746 7129 2748
rect 7153 2746 7209 2748
rect 7233 2746 7289 2748
rect 6993 2694 7039 2746
rect 7039 2694 7049 2746
rect 7073 2694 7103 2746
rect 7103 2694 7115 2746
rect 7115 2694 7129 2746
rect 7153 2694 7167 2746
rect 7167 2694 7179 2746
rect 7179 2694 7209 2746
rect 7233 2694 7243 2746
rect 7243 2694 7289 2746
rect 6993 2692 7049 2694
rect 7073 2692 7129 2694
rect 7153 2692 7209 2694
rect 7233 2692 7289 2694
rect 10874 10376 10930 10432
rect 9408 10362 9464 10364
rect 9488 10362 9544 10364
rect 9568 10362 9624 10364
rect 9648 10362 9704 10364
rect 9408 10310 9454 10362
rect 9454 10310 9464 10362
rect 9488 10310 9518 10362
rect 9518 10310 9530 10362
rect 9530 10310 9544 10362
rect 9568 10310 9582 10362
rect 9582 10310 9594 10362
rect 9594 10310 9624 10362
rect 9648 10310 9658 10362
rect 9658 10310 9704 10362
rect 9408 10308 9464 10310
rect 9488 10308 9544 10310
rect 9568 10308 9624 10310
rect 9648 10308 9704 10310
rect 10068 9818 10124 9820
rect 10148 9818 10204 9820
rect 10228 9818 10284 9820
rect 10308 9818 10364 9820
rect 10068 9766 10114 9818
rect 10114 9766 10124 9818
rect 10148 9766 10178 9818
rect 10178 9766 10190 9818
rect 10190 9766 10204 9818
rect 10228 9766 10242 9818
rect 10242 9766 10254 9818
rect 10254 9766 10284 9818
rect 10308 9766 10318 9818
rect 10318 9766 10364 9818
rect 10068 9764 10124 9766
rect 10148 9764 10204 9766
rect 10228 9764 10284 9766
rect 10308 9764 10364 9766
rect 9408 9274 9464 9276
rect 9488 9274 9544 9276
rect 9568 9274 9624 9276
rect 9648 9274 9704 9276
rect 9408 9222 9454 9274
rect 9454 9222 9464 9274
rect 9488 9222 9518 9274
rect 9518 9222 9530 9274
rect 9530 9222 9544 9274
rect 9568 9222 9582 9274
rect 9582 9222 9594 9274
rect 9594 9222 9624 9274
rect 9648 9222 9658 9274
rect 9658 9222 9704 9274
rect 9408 9220 9464 9222
rect 9488 9220 9544 9222
rect 9568 9220 9624 9222
rect 9648 9220 9704 9222
rect 9408 8186 9464 8188
rect 9488 8186 9544 8188
rect 9568 8186 9624 8188
rect 9648 8186 9704 8188
rect 9408 8134 9454 8186
rect 9454 8134 9464 8186
rect 9488 8134 9518 8186
rect 9518 8134 9530 8186
rect 9530 8134 9544 8186
rect 9568 8134 9582 8186
rect 9582 8134 9594 8186
rect 9594 8134 9624 8186
rect 9648 8134 9658 8186
rect 9658 8134 9704 8186
rect 9408 8132 9464 8134
rect 9488 8132 9544 8134
rect 9568 8132 9624 8134
rect 9648 8132 9704 8134
rect 10068 8730 10124 8732
rect 10148 8730 10204 8732
rect 10228 8730 10284 8732
rect 10308 8730 10364 8732
rect 10068 8678 10114 8730
rect 10114 8678 10124 8730
rect 10148 8678 10178 8730
rect 10178 8678 10190 8730
rect 10190 8678 10204 8730
rect 10228 8678 10242 8730
rect 10242 8678 10254 8730
rect 10254 8678 10284 8730
rect 10308 8678 10318 8730
rect 10318 8678 10364 8730
rect 10068 8676 10124 8678
rect 10148 8676 10204 8678
rect 10228 8676 10284 8678
rect 10308 8676 10364 8678
rect 9408 7098 9464 7100
rect 9488 7098 9544 7100
rect 9568 7098 9624 7100
rect 9648 7098 9704 7100
rect 9408 7046 9454 7098
rect 9454 7046 9464 7098
rect 9488 7046 9518 7098
rect 9518 7046 9530 7098
rect 9530 7046 9544 7098
rect 9568 7046 9582 7098
rect 9582 7046 9594 7098
rect 9594 7046 9624 7098
rect 9648 7046 9658 7098
rect 9658 7046 9704 7098
rect 9408 7044 9464 7046
rect 9488 7044 9544 7046
rect 9568 7044 9624 7046
rect 9648 7044 9704 7046
rect 9408 6010 9464 6012
rect 9488 6010 9544 6012
rect 9568 6010 9624 6012
rect 9648 6010 9704 6012
rect 9408 5958 9454 6010
rect 9454 5958 9464 6010
rect 9488 5958 9518 6010
rect 9518 5958 9530 6010
rect 9530 5958 9544 6010
rect 9568 5958 9582 6010
rect 9582 5958 9594 6010
rect 9594 5958 9624 6010
rect 9648 5958 9658 6010
rect 9658 5958 9704 6010
rect 9408 5956 9464 5958
rect 9488 5956 9544 5958
rect 9568 5956 9624 5958
rect 9648 5956 9704 5958
rect 10068 7642 10124 7644
rect 10148 7642 10204 7644
rect 10228 7642 10284 7644
rect 10308 7642 10364 7644
rect 10068 7590 10114 7642
rect 10114 7590 10124 7642
rect 10148 7590 10178 7642
rect 10178 7590 10190 7642
rect 10190 7590 10204 7642
rect 10228 7590 10242 7642
rect 10242 7590 10254 7642
rect 10254 7590 10284 7642
rect 10308 7590 10318 7642
rect 10318 7590 10364 7642
rect 10068 7588 10124 7590
rect 10148 7588 10204 7590
rect 10228 7588 10284 7590
rect 10308 7588 10364 7590
rect 10068 6554 10124 6556
rect 10148 6554 10204 6556
rect 10228 6554 10284 6556
rect 10308 6554 10364 6556
rect 10068 6502 10114 6554
rect 10114 6502 10124 6554
rect 10148 6502 10178 6554
rect 10178 6502 10190 6554
rect 10190 6502 10204 6554
rect 10228 6502 10242 6554
rect 10242 6502 10254 6554
rect 10254 6502 10284 6554
rect 10308 6502 10318 6554
rect 10318 6502 10364 6554
rect 10068 6500 10124 6502
rect 10148 6500 10204 6502
rect 10228 6500 10284 6502
rect 10308 6500 10364 6502
rect 9408 4922 9464 4924
rect 9488 4922 9544 4924
rect 9568 4922 9624 4924
rect 9648 4922 9704 4924
rect 9408 4870 9454 4922
rect 9454 4870 9464 4922
rect 9488 4870 9518 4922
rect 9518 4870 9530 4922
rect 9530 4870 9544 4922
rect 9568 4870 9582 4922
rect 9582 4870 9594 4922
rect 9594 4870 9624 4922
rect 9648 4870 9658 4922
rect 9658 4870 9704 4922
rect 9408 4868 9464 4870
rect 9488 4868 9544 4870
rect 9568 4868 9624 4870
rect 9648 4868 9704 4870
rect 10068 5466 10124 5468
rect 10148 5466 10204 5468
rect 10228 5466 10284 5468
rect 10308 5466 10364 5468
rect 10068 5414 10114 5466
rect 10114 5414 10124 5466
rect 10148 5414 10178 5466
rect 10178 5414 10190 5466
rect 10190 5414 10204 5466
rect 10228 5414 10242 5466
rect 10242 5414 10254 5466
rect 10254 5414 10284 5466
rect 10308 5414 10318 5466
rect 10318 5414 10364 5466
rect 10068 5412 10124 5414
rect 10148 5412 10204 5414
rect 10228 5412 10284 5414
rect 10308 5412 10364 5414
rect 10068 4378 10124 4380
rect 10148 4378 10204 4380
rect 10228 4378 10284 4380
rect 10308 4378 10364 4380
rect 10068 4326 10114 4378
rect 10114 4326 10124 4378
rect 10148 4326 10178 4378
rect 10178 4326 10190 4378
rect 10190 4326 10204 4378
rect 10228 4326 10242 4378
rect 10242 4326 10254 4378
rect 10254 4326 10284 4378
rect 10308 4326 10318 4378
rect 10318 4326 10364 4378
rect 10068 4324 10124 4326
rect 10148 4324 10204 4326
rect 10228 4324 10284 4326
rect 10308 4324 10364 4326
rect 9408 3834 9464 3836
rect 9488 3834 9544 3836
rect 9568 3834 9624 3836
rect 9648 3834 9704 3836
rect 9408 3782 9454 3834
rect 9454 3782 9464 3834
rect 9488 3782 9518 3834
rect 9518 3782 9530 3834
rect 9530 3782 9544 3834
rect 9568 3782 9582 3834
rect 9582 3782 9594 3834
rect 9594 3782 9624 3834
rect 9648 3782 9658 3834
rect 9658 3782 9704 3834
rect 9408 3780 9464 3782
rect 9488 3780 9544 3782
rect 9568 3780 9624 3782
rect 9648 3780 9704 3782
rect 10068 3290 10124 3292
rect 10148 3290 10204 3292
rect 10228 3290 10284 3292
rect 10308 3290 10364 3292
rect 10068 3238 10114 3290
rect 10114 3238 10124 3290
rect 10148 3238 10178 3290
rect 10178 3238 10190 3290
rect 10190 3238 10204 3290
rect 10228 3238 10242 3290
rect 10242 3238 10254 3290
rect 10254 3238 10284 3290
rect 10308 3238 10318 3290
rect 10318 3238 10364 3290
rect 10068 3236 10124 3238
rect 10148 3236 10204 3238
rect 10228 3236 10284 3238
rect 10308 3236 10364 3238
rect 9408 2746 9464 2748
rect 9488 2746 9544 2748
rect 9568 2746 9624 2748
rect 9648 2746 9704 2748
rect 9408 2694 9454 2746
rect 9454 2694 9464 2746
rect 9488 2694 9518 2746
rect 9518 2694 9530 2746
rect 9530 2694 9544 2746
rect 9568 2694 9582 2746
rect 9582 2694 9594 2746
rect 9594 2694 9624 2746
rect 9648 2694 9658 2746
rect 9658 2694 9704 2746
rect 9408 2692 9464 2694
rect 9488 2692 9544 2694
rect 9568 2692 9624 2694
rect 9648 2692 9704 2694
rect 10874 3304 10930 3360
rect 5238 2202 5294 2204
rect 5318 2202 5374 2204
rect 5398 2202 5454 2204
rect 5478 2202 5534 2204
rect 5238 2150 5284 2202
rect 5284 2150 5294 2202
rect 5318 2150 5348 2202
rect 5348 2150 5360 2202
rect 5360 2150 5374 2202
rect 5398 2150 5412 2202
rect 5412 2150 5424 2202
rect 5424 2150 5454 2202
rect 5478 2150 5488 2202
rect 5488 2150 5534 2202
rect 5238 2148 5294 2150
rect 5318 2148 5374 2150
rect 5398 2148 5454 2150
rect 5478 2148 5534 2150
rect 7653 2202 7709 2204
rect 7733 2202 7789 2204
rect 7813 2202 7869 2204
rect 7893 2202 7949 2204
rect 7653 2150 7699 2202
rect 7699 2150 7709 2202
rect 7733 2150 7763 2202
rect 7763 2150 7775 2202
rect 7775 2150 7789 2202
rect 7813 2150 7827 2202
rect 7827 2150 7839 2202
rect 7839 2150 7869 2202
rect 7893 2150 7903 2202
rect 7903 2150 7949 2202
rect 7653 2148 7709 2150
rect 7733 2148 7789 2150
rect 7813 2148 7869 2150
rect 7893 2148 7949 2150
rect 10068 2202 10124 2204
rect 10148 2202 10204 2204
rect 10228 2202 10284 2204
rect 10308 2202 10364 2204
rect 10068 2150 10114 2202
rect 10114 2150 10124 2202
rect 10148 2150 10178 2202
rect 10178 2150 10190 2202
rect 10190 2150 10204 2202
rect 10228 2150 10242 2202
rect 10242 2150 10254 2202
rect 10254 2150 10284 2202
rect 10308 2150 10318 2202
rect 10318 2150 10364 2202
rect 10068 2148 10124 2150
rect 10148 2148 10204 2150
rect 10228 2148 10284 2150
rect 10308 2148 10364 2150
<< metal3 >>
rect 2153 11456 2469 11457
rect 2153 11392 2159 11456
rect 2223 11392 2239 11456
rect 2303 11392 2319 11456
rect 2383 11392 2399 11456
rect 2463 11392 2469 11456
rect 2153 11391 2469 11392
rect 4568 11456 4884 11457
rect 4568 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4814 11456
rect 4878 11392 4884 11456
rect 4568 11391 4884 11392
rect 6983 11456 7299 11457
rect 6983 11392 6989 11456
rect 7053 11392 7069 11456
rect 7133 11392 7149 11456
rect 7213 11392 7229 11456
rect 7293 11392 7299 11456
rect 6983 11391 7299 11392
rect 9398 11456 9714 11457
rect 9398 11392 9404 11456
rect 9468 11392 9484 11456
rect 9548 11392 9564 11456
rect 9628 11392 9644 11456
rect 9708 11392 9714 11456
rect 9398 11391 9714 11392
rect 2813 10912 3129 10913
rect 2813 10848 2819 10912
rect 2883 10848 2899 10912
rect 2963 10848 2979 10912
rect 3043 10848 3059 10912
rect 3123 10848 3129 10912
rect 2813 10847 3129 10848
rect 5228 10912 5544 10913
rect 5228 10848 5234 10912
rect 5298 10848 5314 10912
rect 5378 10848 5394 10912
rect 5458 10848 5474 10912
rect 5538 10848 5544 10912
rect 5228 10847 5544 10848
rect 7643 10912 7959 10913
rect 7643 10848 7649 10912
rect 7713 10848 7729 10912
rect 7793 10848 7809 10912
rect 7873 10848 7889 10912
rect 7953 10848 7959 10912
rect 7643 10847 7959 10848
rect 10058 10912 10374 10913
rect 10058 10848 10064 10912
rect 10128 10848 10144 10912
rect 10208 10848 10224 10912
rect 10288 10848 10304 10912
rect 10368 10848 10374 10912
rect 10058 10847 10374 10848
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 10869 10434 10935 10437
rect 11154 10434 11954 10464
rect 10869 10432 11954 10434
rect 10869 10376 10874 10432
rect 10930 10376 11954 10432
rect 10869 10374 11954 10376
rect 10869 10371 10935 10374
rect 2153 10368 2469 10369
rect 2153 10304 2159 10368
rect 2223 10304 2239 10368
rect 2303 10304 2319 10368
rect 2383 10304 2399 10368
rect 2463 10304 2469 10368
rect 2153 10303 2469 10304
rect 4568 10368 4884 10369
rect 4568 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4734 10368
rect 4798 10304 4814 10368
rect 4878 10304 4884 10368
rect 4568 10303 4884 10304
rect 6983 10368 7299 10369
rect 6983 10304 6989 10368
rect 7053 10304 7069 10368
rect 7133 10304 7149 10368
rect 7213 10304 7229 10368
rect 7293 10304 7299 10368
rect 6983 10303 7299 10304
rect 9398 10368 9714 10369
rect 9398 10304 9404 10368
rect 9468 10304 9484 10368
rect 9548 10304 9564 10368
rect 9628 10304 9644 10368
rect 9708 10304 9714 10368
rect 11154 10344 11954 10374
rect 9398 10303 9714 10304
rect 2813 9824 3129 9825
rect 2813 9760 2819 9824
rect 2883 9760 2899 9824
rect 2963 9760 2979 9824
rect 3043 9760 3059 9824
rect 3123 9760 3129 9824
rect 2813 9759 3129 9760
rect 5228 9824 5544 9825
rect 5228 9760 5234 9824
rect 5298 9760 5314 9824
rect 5378 9760 5394 9824
rect 5458 9760 5474 9824
rect 5538 9760 5544 9824
rect 5228 9759 5544 9760
rect 7643 9824 7959 9825
rect 7643 9760 7649 9824
rect 7713 9760 7729 9824
rect 7793 9760 7809 9824
rect 7873 9760 7889 9824
rect 7953 9760 7959 9824
rect 7643 9759 7959 9760
rect 10058 9824 10374 9825
rect 10058 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10374 9824
rect 10058 9759 10374 9760
rect 2153 9280 2469 9281
rect 2153 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2399 9280
rect 2463 9216 2469 9280
rect 2153 9215 2469 9216
rect 4568 9280 4884 9281
rect 4568 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4814 9280
rect 4878 9216 4884 9280
rect 4568 9215 4884 9216
rect 6983 9280 7299 9281
rect 6983 9216 6989 9280
rect 7053 9216 7069 9280
rect 7133 9216 7149 9280
rect 7213 9216 7229 9280
rect 7293 9216 7299 9280
rect 6983 9215 7299 9216
rect 9398 9280 9714 9281
rect 9398 9216 9404 9280
rect 9468 9216 9484 9280
rect 9548 9216 9564 9280
rect 9628 9216 9644 9280
rect 9708 9216 9714 9280
rect 9398 9215 9714 9216
rect 2813 8736 3129 8737
rect 2813 8672 2819 8736
rect 2883 8672 2899 8736
rect 2963 8672 2979 8736
rect 3043 8672 3059 8736
rect 3123 8672 3129 8736
rect 2813 8671 3129 8672
rect 5228 8736 5544 8737
rect 5228 8672 5234 8736
rect 5298 8672 5314 8736
rect 5378 8672 5394 8736
rect 5458 8672 5474 8736
rect 5538 8672 5544 8736
rect 5228 8671 5544 8672
rect 7643 8736 7959 8737
rect 7643 8672 7649 8736
rect 7713 8672 7729 8736
rect 7793 8672 7809 8736
rect 7873 8672 7889 8736
rect 7953 8672 7959 8736
rect 7643 8671 7959 8672
rect 10058 8736 10374 8737
rect 10058 8672 10064 8736
rect 10128 8672 10144 8736
rect 10208 8672 10224 8736
rect 10288 8672 10304 8736
rect 10368 8672 10374 8736
rect 10058 8671 10374 8672
rect 2153 8192 2469 8193
rect 2153 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2399 8192
rect 2463 8128 2469 8192
rect 2153 8127 2469 8128
rect 4568 8192 4884 8193
rect 4568 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4814 8192
rect 4878 8128 4884 8192
rect 4568 8127 4884 8128
rect 6983 8192 7299 8193
rect 6983 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7229 8192
rect 7293 8128 7299 8192
rect 6983 8127 7299 8128
rect 9398 8192 9714 8193
rect 9398 8128 9404 8192
rect 9468 8128 9484 8192
rect 9548 8128 9564 8192
rect 9628 8128 9644 8192
rect 9708 8128 9714 8192
rect 9398 8127 9714 8128
rect 2813 7648 3129 7649
rect 2813 7584 2819 7648
rect 2883 7584 2899 7648
rect 2963 7584 2979 7648
rect 3043 7584 3059 7648
rect 3123 7584 3129 7648
rect 2813 7583 3129 7584
rect 5228 7648 5544 7649
rect 5228 7584 5234 7648
rect 5298 7584 5314 7648
rect 5378 7584 5394 7648
rect 5458 7584 5474 7648
rect 5538 7584 5544 7648
rect 5228 7583 5544 7584
rect 7643 7648 7959 7649
rect 7643 7584 7649 7648
rect 7713 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7889 7648
rect 7953 7584 7959 7648
rect 7643 7583 7959 7584
rect 10058 7648 10374 7649
rect 10058 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10374 7648
rect 10058 7583 10374 7584
rect 2153 7104 2469 7105
rect 2153 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2399 7104
rect 2463 7040 2469 7104
rect 2153 7039 2469 7040
rect 4568 7104 4884 7105
rect 4568 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4814 7104
rect 4878 7040 4884 7104
rect 4568 7039 4884 7040
rect 6983 7104 7299 7105
rect 6983 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7229 7104
rect 7293 7040 7299 7104
rect 6983 7039 7299 7040
rect 9398 7104 9714 7105
rect 9398 7040 9404 7104
rect 9468 7040 9484 7104
rect 9548 7040 9564 7104
rect 9628 7040 9644 7104
rect 9708 7040 9714 7104
rect 9398 7039 9714 7040
rect 2813 6560 3129 6561
rect 2813 6496 2819 6560
rect 2883 6496 2899 6560
rect 2963 6496 2979 6560
rect 3043 6496 3059 6560
rect 3123 6496 3129 6560
rect 2813 6495 3129 6496
rect 5228 6560 5544 6561
rect 5228 6496 5234 6560
rect 5298 6496 5314 6560
rect 5378 6496 5394 6560
rect 5458 6496 5474 6560
rect 5538 6496 5544 6560
rect 5228 6495 5544 6496
rect 7643 6560 7959 6561
rect 7643 6496 7649 6560
rect 7713 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7889 6560
rect 7953 6496 7959 6560
rect 7643 6495 7959 6496
rect 10058 6560 10374 6561
rect 10058 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10374 6560
rect 10058 6495 10374 6496
rect 2153 6016 2469 6017
rect 2153 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2399 6016
rect 2463 5952 2469 6016
rect 2153 5951 2469 5952
rect 4568 6016 4884 6017
rect 4568 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4814 6016
rect 4878 5952 4884 6016
rect 4568 5951 4884 5952
rect 6983 6016 7299 6017
rect 6983 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7229 6016
rect 7293 5952 7299 6016
rect 6983 5951 7299 5952
rect 9398 6016 9714 6017
rect 9398 5952 9404 6016
rect 9468 5952 9484 6016
rect 9548 5952 9564 6016
rect 9628 5952 9644 6016
rect 9708 5952 9714 6016
rect 9398 5951 9714 5952
rect 2813 5472 3129 5473
rect 2813 5408 2819 5472
rect 2883 5408 2899 5472
rect 2963 5408 2979 5472
rect 3043 5408 3059 5472
rect 3123 5408 3129 5472
rect 2813 5407 3129 5408
rect 5228 5472 5544 5473
rect 5228 5408 5234 5472
rect 5298 5408 5314 5472
rect 5378 5408 5394 5472
rect 5458 5408 5474 5472
rect 5538 5408 5544 5472
rect 5228 5407 5544 5408
rect 7643 5472 7959 5473
rect 7643 5408 7649 5472
rect 7713 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7889 5472
rect 7953 5408 7959 5472
rect 7643 5407 7959 5408
rect 10058 5472 10374 5473
rect 10058 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10374 5472
rect 10058 5407 10374 5408
rect 2153 4928 2469 4929
rect 2153 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2399 4928
rect 2463 4864 2469 4928
rect 2153 4863 2469 4864
rect 4568 4928 4884 4929
rect 4568 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4814 4928
rect 4878 4864 4884 4928
rect 4568 4863 4884 4864
rect 6983 4928 7299 4929
rect 6983 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7229 4928
rect 7293 4864 7299 4928
rect 6983 4863 7299 4864
rect 9398 4928 9714 4929
rect 9398 4864 9404 4928
rect 9468 4864 9484 4928
rect 9548 4864 9564 4928
rect 9628 4864 9644 4928
rect 9708 4864 9714 4928
rect 9398 4863 9714 4864
rect 2813 4384 3129 4385
rect 2813 4320 2819 4384
rect 2883 4320 2899 4384
rect 2963 4320 2979 4384
rect 3043 4320 3059 4384
rect 3123 4320 3129 4384
rect 2813 4319 3129 4320
rect 5228 4384 5544 4385
rect 5228 4320 5234 4384
rect 5298 4320 5314 4384
rect 5378 4320 5394 4384
rect 5458 4320 5474 4384
rect 5538 4320 5544 4384
rect 5228 4319 5544 4320
rect 7643 4384 7959 4385
rect 7643 4320 7649 4384
rect 7713 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7889 4384
rect 7953 4320 7959 4384
rect 7643 4319 7959 4320
rect 10058 4384 10374 4385
rect 10058 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10374 4384
rect 10058 4319 10374 4320
rect 2153 3840 2469 3841
rect 2153 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2399 3840
rect 2463 3776 2469 3840
rect 2153 3775 2469 3776
rect 4568 3840 4884 3841
rect 4568 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4814 3840
rect 4878 3776 4884 3840
rect 4568 3775 4884 3776
rect 6983 3840 7299 3841
rect 6983 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7229 3840
rect 7293 3776 7299 3840
rect 6983 3775 7299 3776
rect 9398 3840 9714 3841
rect 9398 3776 9404 3840
rect 9468 3776 9484 3840
rect 9548 3776 9564 3840
rect 9628 3776 9644 3840
rect 9708 3776 9714 3840
rect 9398 3775 9714 3776
rect 4061 3498 4127 3501
rect 2638 3496 4127 3498
rect 2638 3440 4066 3496
rect 4122 3440 4127 3496
rect 2638 3438 4127 3440
rect 0 3362 800 3392
rect 2638 3362 2698 3438
rect 4061 3435 4127 3438
rect 0 3302 2698 3362
rect 10869 3362 10935 3365
rect 11154 3362 11954 3392
rect 10869 3360 11954 3362
rect 10869 3304 10874 3360
rect 10930 3304 11954 3360
rect 10869 3302 11954 3304
rect 0 3272 800 3302
rect 10869 3299 10935 3302
rect 2813 3296 3129 3297
rect 2813 3232 2819 3296
rect 2883 3232 2899 3296
rect 2963 3232 2979 3296
rect 3043 3232 3059 3296
rect 3123 3232 3129 3296
rect 2813 3231 3129 3232
rect 5228 3296 5544 3297
rect 5228 3232 5234 3296
rect 5298 3232 5314 3296
rect 5378 3232 5394 3296
rect 5458 3232 5474 3296
rect 5538 3232 5544 3296
rect 5228 3231 5544 3232
rect 7643 3296 7959 3297
rect 7643 3232 7649 3296
rect 7713 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7889 3296
rect 7953 3232 7959 3296
rect 7643 3231 7959 3232
rect 10058 3296 10374 3297
rect 10058 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10374 3296
rect 11154 3272 11954 3302
rect 10058 3231 10374 3232
rect 2153 2752 2469 2753
rect 2153 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2399 2752
rect 2463 2688 2469 2752
rect 2153 2687 2469 2688
rect 4568 2752 4884 2753
rect 4568 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4814 2752
rect 4878 2688 4884 2752
rect 4568 2687 4884 2688
rect 6983 2752 7299 2753
rect 6983 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7229 2752
rect 7293 2688 7299 2752
rect 6983 2687 7299 2688
rect 9398 2752 9714 2753
rect 9398 2688 9404 2752
rect 9468 2688 9484 2752
rect 9548 2688 9564 2752
rect 9628 2688 9644 2752
rect 9708 2688 9714 2752
rect 9398 2687 9714 2688
rect 2813 2208 3129 2209
rect 2813 2144 2819 2208
rect 2883 2144 2899 2208
rect 2963 2144 2979 2208
rect 3043 2144 3059 2208
rect 3123 2144 3129 2208
rect 2813 2143 3129 2144
rect 5228 2208 5544 2209
rect 5228 2144 5234 2208
rect 5298 2144 5314 2208
rect 5378 2144 5394 2208
rect 5458 2144 5474 2208
rect 5538 2144 5544 2208
rect 5228 2143 5544 2144
rect 7643 2208 7959 2209
rect 7643 2144 7649 2208
rect 7713 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7889 2208
rect 7953 2144 7959 2208
rect 7643 2143 7959 2144
rect 10058 2208 10374 2209
rect 10058 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10374 2208
rect 10058 2143 10374 2144
<< via3 >>
rect 2159 11452 2223 11456
rect 2159 11396 2163 11452
rect 2163 11396 2219 11452
rect 2219 11396 2223 11452
rect 2159 11392 2223 11396
rect 2239 11452 2303 11456
rect 2239 11396 2243 11452
rect 2243 11396 2299 11452
rect 2299 11396 2303 11452
rect 2239 11392 2303 11396
rect 2319 11452 2383 11456
rect 2319 11396 2323 11452
rect 2323 11396 2379 11452
rect 2379 11396 2383 11452
rect 2319 11392 2383 11396
rect 2399 11452 2463 11456
rect 2399 11396 2403 11452
rect 2403 11396 2459 11452
rect 2459 11396 2463 11452
rect 2399 11392 2463 11396
rect 4574 11452 4638 11456
rect 4574 11396 4578 11452
rect 4578 11396 4634 11452
rect 4634 11396 4638 11452
rect 4574 11392 4638 11396
rect 4654 11452 4718 11456
rect 4654 11396 4658 11452
rect 4658 11396 4714 11452
rect 4714 11396 4718 11452
rect 4654 11392 4718 11396
rect 4734 11452 4798 11456
rect 4734 11396 4738 11452
rect 4738 11396 4794 11452
rect 4794 11396 4798 11452
rect 4734 11392 4798 11396
rect 4814 11452 4878 11456
rect 4814 11396 4818 11452
rect 4818 11396 4874 11452
rect 4874 11396 4878 11452
rect 4814 11392 4878 11396
rect 6989 11452 7053 11456
rect 6989 11396 6993 11452
rect 6993 11396 7049 11452
rect 7049 11396 7053 11452
rect 6989 11392 7053 11396
rect 7069 11452 7133 11456
rect 7069 11396 7073 11452
rect 7073 11396 7129 11452
rect 7129 11396 7133 11452
rect 7069 11392 7133 11396
rect 7149 11452 7213 11456
rect 7149 11396 7153 11452
rect 7153 11396 7209 11452
rect 7209 11396 7213 11452
rect 7149 11392 7213 11396
rect 7229 11452 7293 11456
rect 7229 11396 7233 11452
rect 7233 11396 7289 11452
rect 7289 11396 7293 11452
rect 7229 11392 7293 11396
rect 9404 11452 9468 11456
rect 9404 11396 9408 11452
rect 9408 11396 9464 11452
rect 9464 11396 9468 11452
rect 9404 11392 9468 11396
rect 9484 11452 9548 11456
rect 9484 11396 9488 11452
rect 9488 11396 9544 11452
rect 9544 11396 9548 11452
rect 9484 11392 9548 11396
rect 9564 11452 9628 11456
rect 9564 11396 9568 11452
rect 9568 11396 9624 11452
rect 9624 11396 9628 11452
rect 9564 11392 9628 11396
rect 9644 11452 9708 11456
rect 9644 11396 9648 11452
rect 9648 11396 9704 11452
rect 9704 11396 9708 11452
rect 9644 11392 9708 11396
rect 2819 10908 2883 10912
rect 2819 10852 2823 10908
rect 2823 10852 2879 10908
rect 2879 10852 2883 10908
rect 2819 10848 2883 10852
rect 2899 10908 2963 10912
rect 2899 10852 2903 10908
rect 2903 10852 2959 10908
rect 2959 10852 2963 10908
rect 2899 10848 2963 10852
rect 2979 10908 3043 10912
rect 2979 10852 2983 10908
rect 2983 10852 3039 10908
rect 3039 10852 3043 10908
rect 2979 10848 3043 10852
rect 3059 10908 3123 10912
rect 3059 10852 3063 10908
rect 3063 10852 3119 10908
rect 3119 10852 3123 10908
rect 3059 10848 3123 10852
rect 5234 10908 5298 10912
rect 5234 10852 5238 10908
rect 5238 10852 5294 10908
rect 5294 10852 5298 10908
rect 5234 10848 5298 10852
rect 5314 10908 5378 10912
rect 5314 10852 5318 10908
rect 5318 10852 5374 10908
rect 5374 10852 5378 10908
rect 5314 10848 5378 10852
rect 5394 10908 5458 10912
rect 5394 10852 5398 10908
rect 5398 10852 5454 10908
rect 5454 10852 5458 10908
rect 5394 10848 5458 10852
rect 5474 10908 5538 10912
rect 5474 10852 5478 10908
rect 5478 10852 5534 10908
rect 5534 10852 5538 10908
rect 5474 10848 5538 10852
rect 7649 10908 7713 10912
rect 7649 10852 7653 10908
rect 7653 10852 7709 10908
rect 7709 10852 7713 10908
rect 7649 10848 7713 10852
rect 7729 10908 7793 10912
rect 7729 10852 7733 10908
rect 7733 10852 7789 10908
rect 7789 10852 7793 10908
rect 7729 10848 7793 10852
rect 7809 10908 7873 10912
rect 7809 10852 7813 10908
rect 7813 10852 7869 10908
rect 7869 10852 7873 10908
rect 7809 10848 7873 10852
rect 7889 10908 7953 10912
rect 7889 10852 7893 10908
rect 7893 10852 7949 10908
rect 7949 10852 7953 10908
rect 7889 10848 7953 10852
rect 10064 10908 10128 10912
rect 10064 10852 10068 10908
rect 10068 10852 10124 10908
rect 10124 10852 10128 10908
rect 10064 10848 10128 10852
rect 10144 10908 10208 10912
rect 10144 10852 10148 10908
rect 10148 10852 10204 10908
rect 10204 10852 10208 10908
rect 10144 10848 10208 10852
rect 10224 10908 10288 10912
rect 10224 10852 10228 10908
rect 10228 10852 10284 10908
rect 10284 10852 10288 10908
rect 10224 10848 10288 10852
rect 10304 10908 10368 10912
rect 10304 10852 10308 10908
rect 10308 10852 10364 10908
rect 10364 10852 10368 10908
rect 10304 10848 10368 10852
rect 2159 10364 2223 10368
rect 2159 10308 2163 10364
rect 2163 10308 2219 10364
rect 2219 10308 2223 10364
rect 2159 10304 2223 10308
rect 2239 10364 2303 10368
rect 2239 10308 2243 10364
rect 2243 10308 2299 10364
rect 2299 10308 2303 10364
rect 2239 10304 2303 10308
rect 2319 10364 2383 10368
rect 2319 10308 2323 10364
rect 2323 10308 2379 10364
rect 2379 10308 2383 10364
rect 2319 10304 2383 10308
rect 2399 10364 2463 10368
rect 2399 10308 2403 10364
rect 2403 10308 2459 10364
rect 2459 10308 2463 10364
rect 2399 10304 2463 10308
rect 4574 10364 4638 10368
rect 4574 10308 4578 10364
rect 4578 10308 4634 10364
rect 4634 10308 4638 10364
rect 4574 10304 4638 10308
rect 4654 10364 4718 10368
rect 4654 10308 4658 10364
rect 4658 10308 4714 10364
rect 4714 10308 4718 10364
rect 4654 10304 4718 10308
rect 4734 10364 4798 10368
rect 4734 10308 4738 10364
rect 4738 10308 4794 10364
rect 4794 10308 4798 10364
rect 4734 10304 4798 10308
rect 4814 10364 4878 10368
rect 4814 10308 4818 10364
rect 4818 10308 4874 10364
rect 4874 10308 4878 10364
rect 4814 10304 4878 10308
rect 6989 10364 7053 10368
rect 6989 10308 6993 10364
rect 6993 10308 7049 10364
rect 7049 10308 7053 10364
rect 6989 10304 7053 10308
rect 7069 10364 7133 10368
rect 7069 10308 7073 10364
rect 7073 10308 7129 10364
rect 7129 10308 7133 10364
rect 7069 10304 7133 10308
rect 7149 10364 7213 10368
rect 7149 10308 7153 10364
rect 7153 10308 7209 10364
rect 7209 10308 7213 10364
rect 7149 10304 7213 10308
rect 7229 10364 7293 10368
rect 7229 10308 7233 10364
rect 7233 10308 7289 10364
rect 7289 10308 7293 10364
rect 7229 10304 7293 10308
rect 9404 10364 9468 10368
rect 9404 10308 9408 10364
rect 9408 10308 9464 10364
rect 9464 10308 9468 10364
rect 9404 10304 9468 10308
rect 9484 10364 9548 10368
rect 9484 10308 9488 10364
rect 9488 10308 9544 10364
rect 9544 10308 9548 10364
rect 9484 10304 9548 10308
rect 9564 10364 9628 10368
rect 9564 10308 9568 10364
rect 9568 10308 9624 10364
rect 9624 10308 9628 10364
rect 9564 10304 9628 10308
rect 9644 10364 9708 10368
rect 9644 10308 9648 10364
rect 9648 10308 9704 10364
rect 9704 10308 9708 10364
rect 9644 10304 9708 10308
rect 2819 9820 2883 9824
rect 2819 9764 2823 9820
rect 2823 9764 2879 9820
rect 2879 9764 2883 9820
rect 2819 9760 2883 9764
rect 2899 9820 2963 9824
rect 2899 9764 2903 9820
rect 2903 9764 2959 9820
rect 2959 9764 2963 9820
rect 2899 9760 2963 9764
rect 2979 9820 3043 9824
rect 2979 9764 2983 9820
rect 2983 9764 3039 9820
rect 3039 9764 3043 9820
rect 2979 9760 3043 9764
rect 3059 9820 3123 9824
rect 3059 9764 3063 9820
rect 3063 9764 3119 9820
rect 3119 9764 3123 9820
rect 3059 9760 3123 9764
rect 5234 9820 5298 9824
rect 5234 9764 5238 9820
rect 5238 9764 5294 9820
rect 5294 9764 5298 9820
rect 5234 9760 5298 9764
rect 5314 9820 5378 9824
rect 5314 9764 5318 9820
rect 5318 9764 5374 9820
rect 5374 9764 5378 9820
rect 5314 9760 5378 9764
rect 5394 9820 5458 9824
rect 5394 9764 5398 9820
rect 5398 9764 5454 9820
rect 5454 9764 5458 9820
rect 5394 9760 5458 9764
rect 5474 9820 5538 9824
rect 5474 9764 5478 9820
rect 5478 9764 5534 9820
rect 5534 9764 5538 9820
rect 5474 9760 5538 9764
rect 7649 9820 7713 9824
rect 7649 9764 7653 9820
rect 7653 9764 7709 9820
rect 7709 9764 7713 9820
rect 7649 9760 7713 9764
rect 7729 9820 7793 9824
rect 7729 9764 7733 9820
rect 7733 9764 7789 9820
rect 7789 9764 7793 9820
rect 7729 9760 7793 9764
rect 7809 9820 7873 9824
rect 7809 9764 7813 9820
rect 7813 9764 7869 9820
rect 7869 9764 7873 9820
rect 7809 9760 7873 9764
rect 7889 9820 7953 9824
rect 7889 9764 7893 9820
rect 7893 9764 7949 9820
rect 7949 9764 7953 9820
rect 7889 9760 7953 9764
rect 10064 9820 10128 9824
rect 10064 9764 10068 9820
rect 10068 9764 10124 9820
rect 10124 9764 10128 9820
rect 10064 9760 10128 9764
rect 10144 9820 10208 9824
rect 10144 9764 10148 9820
rect 10148 9764 10204 9820
rect 10204 9764 10208 9820
rect 10144 9760 10208 9764
rect 10224 9820 10288 9824
rect 10224 9764 10228 9820
rect 10228 9764 10284 9820
rect 10284 9764 10288 9820
rect 10224 9760 10288 9764
rect 10304 9820 10368 9824
rect 10304 9764 10308 9820
rect 10308 9764 10364 9820
rect 10364 9764 10368 9820
rect 10304 9760 10368 9764
rect 2159 9276 2223 9280
rect 2159 9220 2163 9276
rect 2163 9220 2219 9276
rect 2219 9220 2223 9276
rect 2159 9216 2223 9220
rect 2239 9276 2303 9280
rect 2239 9220 2243 9276
rect 2243 9220 2299 9276
rect 2299 9220 2303 9276
rect 2239 9216 2303 9220
rect 2319 9276 2383 9280
rect 2319 9220 2323 9276
rect 2323 9220 2379 9276
rect 2379 9220 2383 9276
rect 2319 9216 2383 9220
rect 2399 9276 2463 9280
rect 2399 9220 2403 9276
rect 2403 9220 2459 9276
rect 2459 9220 2463 9276
rect 2399 9216 2463 9220
rect 4574 9276 4638 9280
rect 4574 9220 4578 9276
rect 4578 9220 4634 9276
rect 4634 9220 4638 9276
rect 4574 9216 4638 9220
rect 4654 9276 4718 9280
rect 4654 9220 4658 9276
rect 4658 9220 4714 9276
rect 4714 9220 4718 9276
rect 4654 9216 4718 9220
rect 4734 9276 4798 9280
rect 4734 9220 4738 9276
rect 4738 9220 4794 9276
rect 4794 9220 4798 9276
rect 4734 9216 4798 9220
rect 4814 9276 4878 9280
rect 4814 9220 4818 9276
rect 4818 9220 4874 9276
rect 4874 9220 4878 9276
rect 4814 9216 4878 9220
rect 6989 9276 7053 9280
rect 6989 9220 6993 9276
rect 6993 9220 7049 9276
rect 7049 9220 7053 9276
rect 6989 9216 7053 9220
rect 7069 9276 7133 9280
rect 7069 9220 7073 9276
rect 7073 9220 7129 9276
rect 7129 9220 7133 9276
rect 7069 9216 7133 9220
rect 7149 9276 7213 9280
rect 7149 9220 7153 9276
rect 7153 9220 7209 9276
rect 7209 9220 7213 9276
rect 7149 9216 7213 9220
rect 7229 9276 7293 9280
rect 7229 9220 7233 9276
rect 7233 9220 7289 9276
rect 7289 9220 7293 9276
rect 7229 9216 7293 9220
rect 9404 9276 9468 9280
rect 9404 9220 9408 9276
rect 9408 9220 9464 9276
rect 9464 9220 9468 9276
rect 9404 9216 9468 9220
rect 9484 9276 9548 9280
rect 9484 9220 9488 9276
rect 9488 9220 9544 9276
rect 9544 9220 9548 9276
rect 9484 9216 9548 9220
rect 9564 9276 9628 9280
rect 9564 9220 9568 9276
rect 9568 9220 9624 9276
rect 9624 9220 9628 9276
rect 9564 9216 9628 9220
rect 9644 9276 9708 9280
rect 9644 9220 9648 9276
rect 9648 9220 9704 9276
rect 9704 9220 9708 9276
rect 9644 9216 9708 9220
rect 2819 8732 2883 8736
rect 2819 8676 2823 8732
rect 2823 8676 2879 8732
rect 2879 8676 2883 8732
rect 2819 8672 2883 8676
rect 2899 8732 2963 8736
rect 2899 8676 2903 8732
rect 2903 8676 2959 8732
rect 2959 8676 2963 8732
rect 2899 8672 2963 8676
rect 2979 8732 3043 8736
rect 2979 8676 2983 8732
rect 2983 8676 3039 8732
rect 3039 8676 3043 8732
rect 2979 8672 3043 8676
rect 3059 8732 3123 8736
rect 3059 8676 3063 8732
rect 3063 8676 3119 8732
rect 3119 8676 3123 8732
rect 3059 8672 3123 8676
rect 5234 8732 5298 8736
rect 5234 8676 5238 8732
rect 5238 8676 5294 8732
rect 5294 8676 5298 8732
rect 5234 8672 5298 8676
rect 5314 8732 5378 8736
rect 5314 8676 5318 8732
rect 5318 8676 5374 8732
rect 5374 8676 5378 8732
rect 5314 8672 5378 8676
rect 5394 8732 5458 8736
rect 5394 8676 5398 8732
rect 5398 8676 5454 8732
rect 5454 8676 5458 8732
rect 5394 8672 5458 8676
rect 5474 8732 5538 8736
rect 5474 8676 5478 8732
rect 5478 8676 5534 8732
rect 5534 8676 5538 8732
rect 5474 8672 5538 8676
rect 7649 8732 7713 8736
rect 7649 8676 7653 8732
rect 7653 8676 7709 8732
rect 7709 8676 7713 8732
rect 7649 8672 7713 8676
rect 7729 8732 7793 8736
rect 7729 8676 7733 8732
rect 7733 8676 7789 8732
rect 7789 8676 7793 8732
rect 7729 8672 7793 8676
rect 7809 8732 7873 8736
rect 7809 8676 7813 8732
rect 7813 8676 7869 8732
rect 7869 8676 7873 8732
rect 7809 8672 7873 8676
rect 7889 8732 7953 8736
rect 7889 8676 7893 8732
rect 7893 8676 7949 8732
rect 7949 8676 7953 8732
rect 7889 8672 7953 8676
rect 10064 8732 10128 8736
rect 10064 8676 10068 8732
rect 10068 8676 10124 8732
rect 10124 8676 10128 8732
rect 10064 8672 10128 8676
rect 10144 8732 10208 8736
rect 10144 8676 10148 8732
rect 10148 8676 10204 8732
rect 10204 8676 10208 8732
rect 10144 8672 10208 8676
rect 10224 8732 10288 8736
rect 10224 8676 10228 8732
rect 10228 8676 10284 8732
rect 10284 8676 10288 8732
rect 10224 8672 10288 8676
rect 10304 8732 10368 8736
rect 10304 8676 10308 8732
rect 10308 8676 10364 8732
rect 10364 8676 10368 8732
rect 10304 8672 10368 8676
rect 2159 8188 2223 8192
rect 2159 8132 2163 8188
rect 2163 8132 2219 8188
rect 2219 8132 2223 8188
rect 2159 8128 2223 8132
rect 2239 8188 2303 8192
rect 2239 8132 2243 8188
rect 2243 8132 2299 8188
rect 2299 8132 2303 8188
rect 2239 8128 2303 8132
rect 2319 8188 2383 8192
rect 2319 8132 2323 8188
rect 2323 8132 2379 8188
rect 2379 8132 2383 8188
rect 2319 8128 2383 8132
rect 2399 8188 2463 8192
rect 2399 8132 2403 8188
rect 2403 8132 2459 8188
rect 2459 8132 2463 8188
rect 2399 8128 2463 8132
rect 4574 8188 4638 8192
rect 4574 8132 4578 8188
rect 4578 8132 4634 8188
rect 4634 8132 4638 8188
rect 4574 8128 4638 8132
rect 4654 8188 4718 8192
rect 4654 8132 4658 8188
rect 4658 8132 4714 8188
rect 4714 8132 4718 8188
rect 4654 8128 4718 8132
rect 4734 8188 4798 8192
rect 4734 8132 4738 8188
rect 4738 8132 4794 8188
rect 4794 8132 4798 8188
rect 4734 8128 4798 8132
rect 4814 8188 4878 8192
rect 4814 8132 4818 8188
rect 4818 8132 4874 8188
rect 4874 8132 4878 8188
rect 4814 8128 4878 8132
rect 6989 8188 7053 8192
rect 6989 8132 6993 8188
rect 6993 8132 7049 8188
rect 7049 8132 7053 8188
rect 6989 8128 7053 8132
rect 7069 8188 7133 8192
rect 7069 8132 7073 8188
rect 7073 8132 7129 8188
rect 7129 8132 7133 8188
rect 7069 8128 7133 8132
rect 7149 8188 7213 8192
rect 7149 8132 7153 8188
rect 7153 8132 7209 8188
rect 7209 8132 7213 8188
rect 7149 8128 7213 8132
rect 7229 8188 7293 8192
rect 7229 8132 7233 8188
rect 7233 8132 7289 8188
rect 7289 8132 7293 8188
rect 7229 8128 7293 8132
rect 9404 8188 9468 8192
rect 9404 8132 9408 8188
rect 9408 8132 9464 8188
rect 9464 8132 9468 8188
rect 9404 8128 9468 8132
rect 9484 8188 9548 8192
rect 9484 8132 9488 8188
rect 9488 8132 9544 8188
rect 9544 8132 9548 8188
rect 9484 8128 9548 8132
rect 9564 8188 9628 8192
rect 9564 8132 9568 8188
rect 9568 8132 9624 8188
rect 9624 8132 9628 8188
rect 9564 8128 9628 8132
rect 9644 8188 9708 8192
rect 9644 8132 9648 8188
rect 9648 8132 9704 8188
rect 9704 8132 9708 8188
rect 9644 8128 9708 8132
rect 2819 7644 2883 7648
rect 2819 7588 2823 7644
rect 2823 7588 2879 7644
rect 2879 7588 2883 7644
rect 2819 7584 2883 7588
rect 2899 7644 2963 7648
rect 2899 7588 2903 7644
rect 2903 7588 2959 7644
rect 2959 7588 2963 7644
rect 2899 7584 2963 7588
rect 2979 7644 3043 7648
rect 2979 7588 2983 7644
rect 2983 7588 3039 7644
rect 3039 7588 3043 7644
rect 2979 7584 3043 7588
rect 3059 7644 3123 7648
rect 3059 7588 3063 7644
rect 3063 7588 3119 7644
rect 3119 7588 3123 7644
rect 3059 7584 3123 7588
rect 5234 7644 5298 7648
rect 5234 7588 5238 7644
rect 5238 7588 5294 7644
rect 5294 7588 5298 7644
rect 5234 7584 5298 7588
rect 5314 7644 5378 7648
rect 5314 7588 5318 7644
rect 5318 7588 5374 7644
rect 5374 7588 5378 7644
rect 5314 7584 5378 7588
rect 5394 7644 5458 7648
rect 5394 7588 5398 7644
rect 5398 7588 5454 7644
rect 5454 7588 5458 7644
rect 5394 7584 5458 7588
rect 5474 7644 5538 7648
rect 5474 7588 5478 7644
rect 5478 7588 5534 7644
rect 5534 7588 5538 7644
rect 5474 7584 5538 7588
rect 7649 7644 7713 7648
rect 7649 7588 7653 7644
rect 7653 7588 7709 7644
rect 7709 7588 7713 7644
rect 7649 7584 7713 7588
rect 7729 7644 7793 7648
rect 7729 7588 7733 7644
rect 7733 7588 7789 7644
rect 7789 7588 7793 7644
rect 7729 7584 7793 7588
rect 7809 7644 7873 7648
rect 7809 7588 7813 7644
rect 7813 7588 7869 7644
rect 7869 7588 7873 7644
rect 7809 7584 7873 7588
rect 7889 7644 7953 7648
rect 7889 7588 7893 7644
rect 7893 7588 7949 7644
rect 7949 7588 7953 7644
rect 7889 7584 7953 7588
rect 10064 7644 10128 7648
rect 10064 7588 10068 7644
rect 10068 7588 10124 7644
rect 10124 7588 10128 7644
rect 10064 7584 10128 7588
rect 10144 7644 10208 7648
rect 10144 7588 10148 7644
rect 10148 7588 10204 7644
rect 10204 7588 10208 7644
rect 10144 7584 10208 7588
rect 10224 7644 10288 7648
rect 10224 7588 10228 7644
rect 10228 7588 10284 7644
rect 10284 7588 10288 7644
rect 10224 7584 10288 7588
rect 10304 7644 10368 7648
rect 10304 7588 10308 7644
rect 10308 7588 10364 7644
rect 10364 7588 10368 7644
rect 10304 7584 10368 7588
rect 2159 7100 2223 7104
rect 2159 7044 2163 7100
rect 2163 7044 2219 7100
rect 2219 7044 2223 7100
rect 2159 7040 2223 7044
rect 2239 7100 2303 7104
rect 2239 7044 2243 7100
rect 2243 7044 2299 7100
rect 2299 7044 2303 7100
rect 2239 7040 2303 7044
rect 2319 7100 2383 7104
rect 2319 7044 2323 7100
rect 2323 7044 2379 7100
rect 2379 7044 2383 7100
rect 2319 7040 2383 7044
rect 2399 7100 2463 7104
rect 2399 7044 2403 7100
rect 2403 7044 2459 7100
rect 2459 7044 2463 7100
rect 2399 7040 2463 7044
rect 4574 7100 4638 7104
rect 4574 7044 4578 7100
rect 4578 7044 4634 7100
rect 4634 7044 4638 7100
rect 4574 7040 4638 7044
rect 4654 7100 4718 7104
rect 4654 7044 4658 7100
rect 4658 7044 4714 7100
rect 4714 7044 4718 7100
rect 4654 7040 4718 7044
rect 4734 7100 4798 7104
rect 4734 7044 4738 7100
rect 4738 7044 4794 7100
rect 4794 7044 4798 7100
rect 4734 7040 4798 7044
rect 4814 7100 4878 7104
rect 4814 7044 4818 7100
rect 4818 7044 4874 7100
rect 4874 7044 4878 7100
rect 4814 7040 4878 7044
rect 6989 7100 7053 7104
rect 6989 7044 6993 7100
rect 6993 7044 7049 7100
rect 7049 7044 7053 7100
rect 6989 7040 7053 7044
rect 7069 7100 7133 7104
rect 7069 7044 7073 7100
rect 7073 7044 7129 7100
rect 7129 7044 7133 7100
rect 7069 7040 7133 7044
rect 7149 7100 7213 7104
rect 7149 7044 7153 7100
rect 7153 7044 7209 7100
rect 7209 7044 7213 7100
rect 7149 7040 7213 7044
rect 7229 7100 7293 7104
rect 7229 7044 7233 7100
rect 7233 7044 7289 7100
rect 7289 7044 7293 7100
rect 7229 7040 7293 7044
rect 9404 7100 9468 7104
rect 9404 7044 9408 7100
rect 9408 7044 9464 7100
rect 9464 7044 9468 7100
rect 9404 7040 9468 7044
rect 9484 7100 9548 7104
rect 9484 7044 9488 7100
rect 9488 7044 9544 7100
rect 9544 7044 9548 7100
rect 9484 7040 9548 7044
rect 9564 7100 9628 7104
rect 9564 7044 9568 7100
rect 9568 7044 9624 7100
rect 9624 7044 9628 7100
rect 9564 7040 9628 7044
rect 9644 7100 9708 7104
rect 9644 7044 9648 7100
rect 9648 7044 9704 7100
rect 9704 7044 9708 7100
rect 9644 7040 9708 7044
rect 2819 6556 2883 6560
rect 2819 6500 2823 6556
rect 2823 6500 2879 6556
rect 2879 6500 2883 6556
rect 2819 6496 2883 6500
rect 2899 6556 2963 6560
rect 2899 6500 2903 6556
rect 2903 6500 2959 6556
rect 2959 6500 2963 6556
rect 2899 6496 2963 6500
rect 2979 6556 3043 6560
rect 2979 6500 2983 6556
rect 2983 6500 3039 6556
rect 3039 6500 3043 6556
rect 2979 6496 3043 6500
rect 3059 6556 3123 6560
rect 3059 6500 3063 6556
rect 3063 6500 3119 6556
rect 3119 6500 3123 6556
rect 3059 6496 3123 6500
rect 5234 6556 5298 6560
rect 5234 6500 5238 6556
rect 5238 6500 5294 6556
rect 5294 6500 5298 6556
rect 5234 6496 5298 6500
rect 5314 6556 5378 6560
rect 5314 6500 5318 6556
rect 5318 6500 5374 6556
rect 5374 6500 5378 6556
rect 5314 6496 5378 6500
rect 5394 6556 5458 6560
rect 5394 6500 5398 6556
rect 5398 6500 5454 6556
rect 5454 6500 5458 6556
rect 5394 6496 5458 6500
rect 5474 6556 5538 6560
rect 5474 6500 5478 6556
rect 5478 6500 5534 6556
rect 5534 6500 5538 6556
rect 5474 6496 5538 6500
rect 7649 6556 7713 6560
rect 7649 6500 7653 6556
rect 7653 6500 7709 6556
rect 7709 6500 7713 6556
rect 7649 6496 7713 6500
rect 7729 6556 7793 6560
rect 7729 6500 7733 6556
rect 7733 6500 7789 6556
rect 7789 6500 7793 6556
rect 7729 6496 7793 6500
rect 7809 6556 7873 6560
rect 7809 6500 7813 6556
rect 7813 6500 7869 6556
rect 7869 6500 7873 6556
rect 7809 6496 7873 6500
rect 7889 6556 7953 6560
rect 7889 6500 7893 6556
rect 7893 6500 7949 6556
rect 7949 6500 7953 6556
rect 7889 6496 7953 6500
rect 10064 6556 10128 6560
rect 10064 6500 10068 6556
rect 10068 6500 10124 6556
rect 10124 6500 10128 6556
rect 10064 6496 10128 6500
rect 10144 6556 10208 6560
rect 10144 6500 10148 6556
rect 10148 6500 10204 6556
rect 10204 6500 10208 6556
rect 10144 6496 10208 6500
rect 10224 6556 10288 6560
rect 10224 6500 10228 6556
rect 10228 6500 10284 6556
rect 10284 6500 10288 6556
rect 10224 6496 10288 6500
rect 10304 6556 10368 6560
rect 10304 6500 10308 6556
rect 10308 6500 10364 6556
rect 10364 6500 10368 6556
rect 10304 6496 10368 6500
rect 2159 6012 2223 6016
rect 2159 5956 2163 6012
rect 2163 5956 2219 6012
rect 2219 5956 2223 6012
rect 2159 5952 2223 5956
rect 2239 6012 2303 6016
rect 2239 5956 2243 6012
rect 2243 5956 2299 6012
rect 2299 5956 2303 6012
rect 2239 5952 2303 5956
rect 2319 6012 2383 6016
rect 2319 5956 2323 6012
rect 2323 5956 2379 6012
rect 2379 5956 2383 6012
rect 2319 5952 2383 5956
rect 2399 6012 2463 6016
rect 2399 5956 2403 6012
rect 2403 5956 2459 6012
rect 2459 5956 2463 6012
rect 2399 5952 2463 5956
rect 4574 6012 4638 6016
rect 4574 5956 4578 6012
rect 4578 5956 4634 6012
rect 4634 5956 4638 6012
rect 4574 5952 4638 5956
rect 4654 6012 4718 6016
rect 4654 5956 4658 6012
rect 4658 5956 4714 6012
rect 4714 5956 4718 6012
rect 4654 5952 4718 5956
rect 4734 6012 4798 6016
rect 4734 5956 4738 6012
rect 4738 5956 4794 6012
rect 4794 5956 4798 6012
rect 4734 5952 4798 5956
rect 4814 6012 4878 6016
rect 4814 5956 4818 6012
rect 4818 5956 4874 6012
rect 4874 5956 4878 6012
rect 4814 5952 4878 5956
rect 6989 6012 7053 6016
rect 6989 5956 6993 6012
rect 6993 5956 7049 6012
rect 7049 5956 7053 6012
rect 6989 5952 7053 5956
rect 7069 6012 7133 6016
rect 7069 5956 7073 6012
rect 7073 5956 7129 6012
rect 7129 5956 7133 6012
rect 7069 5952 7133 5956
rect 7149 6012 7213 6016
rect 7149 5956 7153 6012
rect 7153 5956 7209 6012
rect 7209 5956 7213 6012
rect 7149 5952 7213 5956
rect 7229 6012 7293 6016
rect 7229 5956 7233 6012
rect 7233 5956 7289 6012
rect 7289 5956 7293 6012
rect 7229 5952 7293 5956
rect 9404 6012 9468 6016
rect 9404 5956 9408 6012
rect 9408 5956 9464 6012
rect 9464 5956 9468 6012
rect 9404 5952 9468 5956
rect 9484 6012 9548 6016
rect 9484 5956 9488 6012
rect 9488 5956 9544 6012
rect 9544 5956 9548 6012
rect 9484 5952 9548 5956
rect 9564 6012 9628 6016
rect 9564 5956 9568 6012
rect 9568 5956 9624 6012
rect 9624 5956 9628 6012
rect 9564 5952 9628 5956
rect 9644 6012 9708 6016
rect 9644 5956 9648 6012
rect 9648 5956 9704 6012
rect 9704 5956 9708 6012
rect 9644 5952 9708 5956
rect 2819 5468 2883 5472
rect 2819 5412 2823 5468
rect 2823 5412 2879 5468
rect 2879 5412 2883 5468
rect 2819 5408 2883 5412
rect 2899 5468 2963 5472
rect 2899 5412 2903 5468
rect 2903 5412 2959 5468
rect 2959 5412 2963 5468
rect 2899 5408 2963 5412
rect 2979 5468 3043 5472
rect 2979 5412 2983 5468
rect 2983 5412 3039 5468
rect 3039 5412 3043 5468
rect 2979 5408 3043 5412
rect 3059 5468 3123 5472
rect 3059 5412 3063 5468
rect 3063 5412 3119 5468
rect 3119 5412 3123 5468
rect 3059 5408 3123 5412
rect 5234 5468 5298 5472
rect 5234 5412 5238 5468
rect 5238 5412 5294 5468
rect 5294 5412 5298 5468
rect 5234 5408 5298 5412
rect 5314 5468 5378 5472
rect 5314 5412 5318 5468
rect 5318 5412 5374 5468
rect 5374 5412 5378 5468
rect 5314 5408 5378 5412
rect 5394 5468 5458 5472
rect 5394 5412 5398 5468
rect 5398 5412 5454 5468
rect 5454 5412 5458 5468
rect 5394 5408 5458 5412
rect 5474 5468 5538 5472
rect 5474 5412 5478 5468
rect 5478 5412 5534 5468
rect 5534 5412 5538 5468
rect 5474 5408 5538 5412
rect 7649 5468 7713 5472
rect 7649 5412 7653 5468
rect 7653 5412 7709 5468
rect 7709 5412 7713 5468
rect 7649 5408 7713 5412
rect 7729 5468 7793 5472
rect 7729 5412 7733 5468
rect 7733 5412 7789 5468
rect 7789 5412 7793 5468
rect 7729 5408 7793 5412
rect 7809 5468 7873 5472
rect 7809 5412 7813 5468
rect 7813 5412 7869 5468
rect 7869 5412 7873 5468
rect 7809 5408 7873 5412
rect 7889 5468 7953 5472
rect 7889 5412 7893 5468
rect 7893 5412 7949 5468
rect 7949 5412 7953 5468
rect 7889 5408 7953 5412
rect 10064 5468 10128 5472
rect 10064 5412 10068 5468
rect 10068 5412 10124 5468
rect 10124 5412 10128 5468
rect 10064 5408 10128 5412
rect 10144 5468 10208 5472
rect 10144 5412 10148 5468
rect 10148 5412 10204 5468
rect 10204 5412 10208 5468
rect 10144 5408 10208 5412
rect 10224 5468 10288 5472
rect 10224 5412 10228 5468
rect 10228 5412 10284 5468
rect 10284 5412 10288 5468
rect 10224 5408 10288 5412
rect 10304 5468 10368 5472
rect 10304 5412 10308 5468
rect 10308 5412 10364 5468
rect 10364 5412 10368 5468
rect 10304 5408 10368 5412
rect 2159 4924 2223 4928
rect 2159 4868 2163 4924
rect 2163 4868 2219 4924
rect 2219 4868 2223 4924
rect 2159 4864 2223 4868
rect 2239 4924 2303 4928
rect 2239 4868 2243 4924
rect 2243 4868 2299 4924
rect 2299 4868 2303 4924
rect 2239 4864 2303 4868
rect 2319 4924 2383 4928
rect 2319 4868 2323 4924
rect 2323 4868 2379 4924
rect 2379 4868 2383 4924
rect 2319 4864 2383 4868
rect 2399 4924 2463 4928
rect 2399 4868 2403 4924
rect 2403 4868 2459 4924
rect 2459 4868 2463 4924
rect 2399 4864 2463 4868
rect 4574 4924 4638 4928
rect 4574 4868 4578 4924
rect 4578 4868 4634 4924
rect 4634 4868 4638 4924
rect 4574 4864 4638 4868
rect 4654 4924 4718 4928
rect 4654 4868 4658 4924
rect 4658 4868 4714 4924
rect 4714 4868 4718 4924
rect 4654 4864 4718 4868
rect 4734 4924 4798 4928
rect 4734 4868 4738 4924
rect 4738 4868 4794 4924
rect 4794 4868 4798 4924
rect 4734 4864 4798 4868
rect 4814 4924 4878 4928
rect 4814 4868 4818 4924
rect 4818 4868 4874 4924
rect 4874 4868 4878 4924
rect 4814 4864 4878 4868
rect 6989 4924 7053 4928
rect 6989 4868 6993 4924
rect 6993 4868 7049 4924
rect 7049 4868 7053 4924
rect 6989 4864 7053 4868
rect 7069 4924 7133 4928
rect 7069 4868 7073 4924
rect 7073 4868 7129 4924
rect 7129 4868 7133 4924
rect 7069 4864 7133 4868
rect 7149 4924 7213 4928
rect 7149 4868 7153 4924
rect 7153 4868 7209 4924
rect 7209 4868 7213 4924
rect 7149 4864 7213 4868
rect 7229 4924 7293 4928
rect 7229 4868 7233 4924
rect 7233 4868 7289 4924
rect 7289 4868 7293 4924
rect 7229 4864 7293 4868
rect 9404 4924 9468 4928
rect 9404 4868 9408 4924
rect 9408 4868 9464 4924
rect 9464 4868 9468 4924
rect 9404 4864 9468 4868
rect 9484 4924 9548 4928
rect 9484 4868 9488 4924
rect 9488 4868 9544 4924
rect 9544 4868 9548 4924
rect 9484 4864 9548 4868
rect 9564 4924 9628 4928
rect 9564 4868 9568 4924
rect 9568 4868 9624 4924
rect 9624 4868 9628 4924
rect 9564 4864 9628 4868
rect 9644 4924 9708 4928
rect 9644 4868 9648 4924
rect 9648 4868 9704 4924
rect 9704 4868 9708 4924
rect 9644 4864 9708 4868
rect 2819 4380 2883 4384
rect 2819 4324 2823 4380
rect 2823 4324 2879 4380
rect 2879 4324 2883 4380
rect 2819 4320 2883 4324
rect 2899 4380 2963 4384
rect 2899 4324 2903 4380
rect 2903 4324 2959 4380
rect 2959 4324 2963 4380
rect 2899 4320 2963 4324
rect 2979 4380 3043 4384
rect 2979 4324 2983 4380
rect 2983 4324 3039 4380
rect 3039 4324 3043 4380
rect 2979 4320 3043 4324
rect 3059 4380 3123 4384
rect 3059 4324 3063 4380
rect 3063 4324 3119 4380
rect 3119 4324 3123 4380
rect 3059 4320 3123 4324
rect 5234 4380 5298 4384
rect 5234 4324 5238 4380
rect 5238 4324 5294 4380
rect 5294 4324 5298 4380
rect 5234 4320 5298 4324
rect 5314 4380 5378 4384
rect 5314 4324 5318 4380
rect 5318 4324 5374 4380
rect 5374 4324 5378 4380
rect 5314 4320 5378 4324
rect 5394 4380 5458 4384
rect 5394 4324 5398 4380
rect 5398 4324 5454 4380
rect 5454 4324 5458 4380
rect 5394 4320 5458 4324
rect 5474 4380 5538 4384
rect 5474 4324 5478 4380
rect 5478 4324 5534 4380
rect 5534 4324 5538 4380
rect 5474 4320 5538 4324
rect 7649 4380 7713 4384
rect 7649 4324 7653 4380
rect 7653 4324 7709 4380
rect 7709 4324 7713 4380
rect 7649 4320 7713 4324
rect 7729 4380 7793 4384
rect 7729 4324 7733 4380
rect 7733 4324 7789 4380
rect 7789 4324 7793 4380
rect 7729 4320 7793 4324
rect 7809 4380 7873 4384
rect 7809 4324 7813 4380
rect 7813 4324 7869 4380
rect 7869 4324 7873 4380
rect 7809 4320 7873 4324
rect 7889 4380 7953 4384
rect 7889 4324 7893 4380
rect 7893 4324 7949 4380
rect 7949 4324 7953 4380
rect 7889 4320 7953 4324
rect 10064 4380 10128 4384
rect 10064 4324 10068 4380
rect 10068 4324 10124 4380
rect 10124 4324 10128 4380
rect 10064 4320 10128 4324
rect 10144 4380 10208 4384
rect 10144 4324 10148 4380
rect 10148 4324 10204 4380
rect 10204 4324 10208 4380
rect 10144 4320 10208 4324
rect 10224 4380 10288 4384
rect 10224 4324 10228 4380
rect 10228 4324 10284 4380
rect 10284 4324 10288 4380
rect 10224 4320 10288 4324
rect 10304 4380 10368 4384
rect 10304 4324 10308 4380
rect 10308 4324 10364 4380
rect 10364 4324 10368 4380
rect 10304 4320 10368 4324
rect 2159 3836 2223 3840
rect 2159 3780 2163 3836
rect 2163 3780 2219 3836
rect 2219 3780 2223 3836
rect 2159 3776 2223 3780
rect 2239 3836 2303 3840
rect 2239 3780 2243 3836
rect 2243 3780 2299 3836
rect 2299 3780 2303 3836
rect 2239 3776 2303 3780
rect 2319 3836 2383 3840
rect 2319 3780 2323 3836
rect 2323 3780 2379 3836
rect 2379 3780 2383 3836
rect 2319 3776 2383 3780
rect 2399 3836 2463 3840
rect 2399 3780 2403 3836
rect 2403 3780 2459 3836
rect 2459 3780 2463 3836
rect 2399 3776 2463 3780
rect 4574 3836 4638 3840
rect 4574 3780 4578 3836
rect 4578 3780 4634 3836
rect 4634 3780 4638 3836
rect 4574 3776 4638 3780
rect 4654 3836 4718 3840
rect 4654 3780 4658 3836
rect 4658 3780 4714 3836
rect 4714 3780 4718 3836
rect 4654 3776 4718 3780
rect 4734 3836 4798 3840
rect 4734 3780 4738 3836
rect 4738 3780 4794 3836
rect 4794 3780 4798 3836
rect 4734 3776 4798 3780
rect 4814 3836 4878 3840
rect 4814 3780 4818 3836
rect 4818 3780 4874 3836
rect 4874 3780 4878 3836
rect 4814 3776 4878 3780
rect 6989 3836 7053 3840
rect 6989 3780 6993 3836
rect 6993 3780 7049 3836
rect 7049 3780 7053 3836
rect 6989 3776 7053 3780
rect 7069 3836 7133 3840
rect 7069 3780 7073 3836
rect 7073 3780 7129 3836
rect 7129 3780 7133 3836
rect 7069 3776 7133 3780
rect 7149 3836 7213 3840
rect 7149 3780 7153 3836
rect 7153 3780 7209 3836
rect 7209 3780 7213 3836
rect 7149 3776 7213 3780
rect 7229 3836 7293 3840
rect 7229 3780 7233 3836
rect 7233 3780 7289 3836
rect 7289 3780 7293 3836
rect 7229 3776 7293 3780
rect 9404 3836 9468 3840
rect 9404 3780 9408 3836
rect 9408 3780 9464 3836
rect 9464 3780 9468 3836
rect 9404 3776 9468 3780
rect 9484 3836 9548 3840
rect 9484 3780 9488 3836
rect 9488 3780 9544 3836
rect 9544 3780 9548 3836
rect 9484 3776 9548 3780
rect 9564 3836 9628 3840
rect 9564 3780 9568 3836
rect 9568 3780 9624 3836
rect 9624 3780 9628 3836
rect 9564 3776 9628 3780
rect 9644 3836 9708 3840
rect 9644 3780 9648 3836
rect 9648 3780 9704 3836
rect 9704 3780 9708 3836
rect 9644 3776 9708 3780
rect 2819 3292 2883 3296
rect 2819 3236 2823 3292
rect 2823 3236 2879 3292
rect 2879 3236 2883 3292
rect 2819 3232 2883 3236
rect 2899 3292 2963 3296
rect 2899 3236 2903 3292
rect 2903 3236 2959 3292
rect 2959 3236 2963 3292
rect 2899 3232 2963 3236
rect 2979 3292 3043 3296
rect 2979 3236 2983 3292
rect 2983 3236 3039 3292
rect 3039 3236 3043 3292
rect 2979 3232 3043 3236
rect 3059 3292 3123 3296
rect 3059 3236 3063 3292
rect 3063 3236 3119 3292
rect 3119 3236 3123 3292
rect 3059 3232 3123 3236
rect 5234 3292 5298 3296
rect 5234 3236 5238 3292
rect 5238 3236 5294 3292
rect 5294 3236 5298 3292
rect 5234 3232 5298 3236
rect 5314 3292 5378 3296
rect 5314 3236 5318 3292
rect 5318 3236 5374 3292
rect 5374 3236 5378 3292
rect 5314 3232 5378 3236
rect 5394 3292 5458 3296
rect 5394 3236 5398 3292
rect 5398 3236 5454 3292
rect 5454 3236 5458 3292
rect 5394 3232 5458 3236
rect 5474 3292 5538 3296
rect 5474 3236 5478 3292
rect 5478 3236 5534 3292
rect 5534 3236 5538 3292
rect 5474 3232 5538 3236
rect 7649 3292 7713 3296
rect 7649 3236 7653 3292
rect 7653 3236 7709 3292
rect 7709 3236 7713 3292
rect 7649 3232 7713 3236
rect 7729 3292 7793 3296
rect 7729 3236 7733 3292
rect 7733 3236 7789 3292
rect 7789 3236 7793 3292
rect 7729 3232 7793 3236
rect 7809 3292 7873 3296
rect 7809 3236 7813 3292
rect 7813 3236 7869 3292
rect 7869 3236 7873 3292
rect 7809 3232 7873 3236
rect 7889 3292 7953 3296
rect 7889 3236 7893 3292
rect 7893 3236 7949 3292
rect 7949 3236 7953 3292
rect 7889 3232 7953 3236
rect 10064 3292 10128 3296
rect 10064 3236 10068 3292
rect 10068 3236 10124 3292
rect 10124 3236 10128 3292
rect 10064 3232 10128 3236
rect 10144 3292 10208 3296
rect 10144 3236 10148 3292
rect 10148 3236 10204 3292
rect 10204 3236 10208 3292
rect 10144 3232 10208 3236
rect 10224 3292 10288 3296
rect 10224 3236 10228 3292
rect 10228 3236 10284 3292
rect 10284 3236 10288 3292
rect 10224 3232 10288 3236
rect 10304 3292 10368 3296
rect 10304 3236 10308 3292
rect 10308 3236 10364 3292
rect 10364 3236 10368 3292
rect 10304 3232 10368 3236
rect 2159 2748 2223 2752
rect 2159 2692 2163 2748
rect 2163 2692 2219 2748
rect 2219 2692 2223 2748
rect 2159 2688 2223 2692
rect 2239 2748 2303 2752
rect 2239 2692 2243 2748
rect 2243 2692 2299 2748
rect 2299 2692 2303 2748
rect 2239 2688 2303 2692
rect 2319 2748 2383 2752
rect 2319 2692 2323 2748
rect 2323 2692 2379 2748
rect 2379 2692 2383 2748
rect 2319 2688 2383 2692
rect 2399 2748 2463 2752
rect 2399 2692 2403 2748
rect 2403 2692 2459 2748
rect 2459 2692 2463 2748
rect 2399 2688 2463 2692
rect 4574 2748 4638 2752
rect 4574 2692 4578 2748
rect 4578 2692 4634 2748
rect 4634 2692 4638 2748
rect 4574 2688 4638 2692
rect 4654 2748 4718 2752
rect 4654 2692 4658 2748
rect 4658 2692 4714 2748
rect 4714 2692 4718 2748
rect 4654 2688 4718 2692
rect 4734 2748 4798 2752
rect 4734 2692 4738 2748
rect 4738 2692 4794 2748
rect 4794 2692 4798 2748
rect 4734 2688 4798 2692
rect 4814 2748 4878 2752
rect 4814 2692 4818 2748
rect 4818 2692 4874 2748
rect 4874 2692 4878 2748
rect 4814 2688 4878 2692
rect 6989 2748 7053 2752
rect 6989 2692 6993 2748
rect 6993 2692 7049 2748
rect 7049 2692 7053 2748
rect 6989 2688 7053 2692
rect 7069 2748 7133 2752
rect 7069 2692 7073 2748
rect 7073 2692 7129 2748
rect 7129 2692 7133 2748
rect 7069 2688 7133 2692
rect 7149 2748 7213 2752
rect 7149 2692 7153 2748
rect 7153 2692 7209 2748
rect 7209 2692 7213 2748
rect 7149 2688 7213 2692
rect 7229 2748 7293 2752
rect 7229 2692 7233 2748
rect 7233 2692 7289 2748
rect 7289 2692 7293 2748
rect 7229 2688 7293 2692
rect 9404 2748 9468 2752
rect 9404 2692 9408 2748
rect 9408 2692 9464 2748
rect 9464 2692 9468 2748
rect 9404 2688 9468 2692
rect 9484 2748 9548 2752
rect 9484 2692 9488 2748
rect 9488 2692 9544 2748
rect 9544 2692 9548 2748
rect 9484 2688 9548 2692
rect 9564 2748 9628 2752
rect 9564 2692 9568 2748
rect 9568 2692 9624 2748
rect 9624 2692 9628 2748
rect 9564 2688 9628 2692
rect 9644 2748 9708 2752
rect 9644 2692 9648 2748
rect 9648 2692 9704 2748
rect 9704 2692 9708 2748
rect 9644 2688 9708 2692
rect 2819 2204 2883 2208
rect 2819 2148 2823 2204
rect 2823 2148 2879 2204
rect 2879 2148 2883 2204
rect 2819 2144 2883 2148
rect 2899 2204 2963 2208
rect 2899 2148 2903 2204
rect 2903 2148 2959 2204
rect 2959 2148 2963 2204
rect 2899 2144 2963 2148
rect 2979 2204 3043 2208
rect 2979 2148 2983 2204
rect 2983 2148 3039 2204
rect 3039 2148 3043 2204
rect 2979 2144 3043 2148
rect 3059 2204 3123 2208
rect 3059 2148 3063 2204
rect 3063 2148 3119 2204
rect 3119 2148 3123 2204
rect 3059 2144 3123 2148
rect 5234 2204 5298 2208
rect 5234 2148 5238 2204
rect 5238 2148 5294 2204
rect 5294 2148 5298 2204
rect 5234 2144 5298 2148
rect 5314 2204 5378 2208
rect 5314 2148 5318 2204
rect 5318 2148 5374 2204
rect 5374 2148 5378 2204
rect 5314 2144 5378 2148
rect 5394 2204 5458 2208
rect 5394 2148 5398 2204
rect 5398 2148 5454 2204
rect 5454 2148 5458 2204
rect 5394 2144 5458 2148
rect 5474 2204 5538 2208
rect 5474 2148 5478 2204
rect 5478 2148 5534 2204
rect 5534 2148 5538 2204
rect 5474 2144 5538 2148
rect 7649 2204 7713 2208
rect 7649 2148 7653 2204
rect 7653 2148 7709 2204
rect 7709 2148 7713 2204
rect 7649 2144 7713 2148
rect 7729 2204 7793 2208
rect 7729 2148 7733 2204
rect 7733 2148 7789 2204
rect 7789 2148 7793 2204
rect 7729 2144 7793 2148
rect 7809 2204 7873 2208
rect 7809 2148 7813 2204
rect 7813 2148 7869 2204
rect 7869 2148 7873 2204
rect 7809 2144 7873 2148
rect 7889 2204 7953 2208
rect 7889 2148 7893 2204
rect 7893 2148 7949 2204
rect 7949 2148 7953 2204
rect 7889 2144 7953 2148
rect 10064 2204 10128 2208
rect 10064 2148 10068 2204
rect 10068 2148 10124 2204
rect 10124 2148 10128 2204
rect 10064 2144 10128 2148
rect 10144 2204 10208 2208
rect 10144 2148 10148 2204
rect 10148 2148 10204 2204
rect 10204 2148 10208 2204
rect 10144 2144 10208 2148
rect 10224 2204 10288 2208
rect 10224 2148 10228 2204
rect 10228 2148 10284 2204
rect 10284 2148 10288 2204
rect 10224 2144 10288 2148
rect 10304 2204 10368 2208
rect 10304 2148 10308 2204
rect 10308 2148 10364 2204
rect 10364 2148 10368 2204
rect 10304 2144 10368 2148
<< metal4 >>
rect 2151 11456 2471 11472
rect 2151 11392 2159 11456
rect 2223 11392 2239 11456
rect 2303 11392 2319 11456
rect 2383 11392 2399 11456
rect 2463 11392 2471 11456
rect 2151 10382 2471 11392
rect 2151 10368 2193 10382
rect 2429 10368 2471 10382
rect 2151 10304 2159 10368
rect 2463 10304 2471 10368
rect 2151 10146 2193 10304
rect 2429 10146 2471 10304
rect 2151 9280 2471 10146
rect 2151 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2399 9280
rect 2463 9216 2471 9280
rect 2151 8192 2471 9216
rect 2151 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2399 8192
rect 2463 8128 2471 8192
rect 2151 8071 2471 8128
rect 2151 7835 2193 8071
rect 2429 7835 2471 8071
rect 2151 7104 2471 7835
rect 2151 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2399 7104
rect 2463 7040 2471 7104
rect 2151 6016 2471 7040
rect 2151 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2399 6016
rect 2463 5952 2471 6016
rect 2151 5760 2471 5952
rect 2151 5524 2193 5760
rect 2429 5524 2471 5760
rect 2151 4928 2471 5524
rect 2151 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2399 4928
rect 2463 4864 2471 4928
rect 2151 3840 2471 4864
rect 2151 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2399 3840
rect 2463 3776 2471 3840
rect 2151 3449 2471 3776
rect 2151 3213 2193 3449
rect 2429 3213 2471 3449
rect 2151 2752 2471 3213
rect 2151 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2399 2752
rect 2463 2688 2471 2752
rect 2151 2128 2471 2688
rect 2811 11042 3131 11472
rect 2811 10912 2853 11042
rect 3089 10912 3131 11042
rect 2811 10848 2819 10912
rect 3123 10848 3131 10912
rect 2811 10806 2853 10848
rect 3089 10806 3131 10848
rect 2811 9824 3131 10806
rect 2811 9760 2819 9824
rect 2883 9760 2899 9824
rect 2963 9760 2979 9824
rect 3043 9760 3059 9824
rect 3123 9760 3131 9824
rect 2811 8736 3131 9760
rect 2811 8672 2819 8736
rect 2883 8731 2899 8736
rect 2963 8731 2979 8736
rect 3043 8731 3059 8736
rect 3123 8672 3131 8736
rect 2811 8495 2853 8672
rect 3089 8495 3131 8672
rect 2811 7648 3131 8495
rect 2811 7584 2819 7648
rect 2883 7584 2899 7648
rect 2963 7584 2979 7648
rect 3043 7584 3059 7648
rect 3123 7584 3131 7648
rect 2811 6560 3131 7584
rect 2811 6496 2819 6560
rect 2883 6496 2899 6560
rect 2963 6496 2979 6560
rect 3043 6496 3059 6560
rect 3123 6496 3131 6560
rect 2811 6420 3131 6496
rect 2811 6184 2853 6420
rect 3089 6184 3131 6420
rect 2811 5472 3131 6184
rect 2811 5408 2819 5472
rect 2883 5408 2899 5472
rect 2963 5408 2979 5472
rect 3043 5408 3059 5472
rect 3123 5408 3131 5472
rect 2811 4384 3131 5408
rect 2811 4320 2819 4384
rect 2883 4320 2899 4384
rect 2963 4320 2979 4384
rect 3043 4320 3059 4384
rect 3123 4320 3131 4384
rect 2811 4109 3131 4320
rect 2811 3873 2853 4109
rect 3089 3873 3131 4109
rect 2811 3296 3131 3873
rect 2811 3232 2819 3296
rect 2883 3232 2899 3296
rect 2963 3232 2979 3296
rect 3043 3232 3059 3296
rect 3123 3232 3131 3296
rect 2811 2208 3131 3232
rect 2811 2144 2819 2208
rect 2883 2144 2899 2208
rect 2963 2144 2979 2208
rect 3043 2144 3059 2208
rect 3123 2144 3131 2208
rect 2811 2128 3131 2144
rect 4566 11456 4886 11472
rect 4566 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4814 11456
rect 4878 11392 4886 11456
rect 4566 10382 4886 11392
rect 4566 10368 4608 10382
rect 4844 10368 4886 10382
rect 4566 10304 4574 10368
rect 4878 10304 4886 10368
rect 4566 10146 4608 10304
rect 4844 10146 4886 10304
rect 4566 9280 4886 10146
rect 4566 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4814 9280
rect 4878 9216 4886 9280
rect 4566 8192 4886 9216
rect 4566 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4814 8192
rect 4878 8128 4886 8192
rect 4566 8071 4886 8128
rect 4566 7835 4608 8071
rect 4844 7835 4886 8071
rect 4566 7104 4886 7835
rect 4566 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4814 7104
rect 4878 7040 4886 7104
rect 4566 6016 4886 7040
rect 4566 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4814 6016
rect 4878 5952 4886 6016
rect 4566 5760 4886 5952
rect 4566 5524 4608 5760
rect 4844 5524 4886 5760
rect 4566 4928 4886 5524
rect 4566 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4814 4928
rect 4878 4864 4886 4928
rect 4566 3840 4886 4864
rect 4566 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4814 3840
rect 4878 3776 4886 3840
rect 4566 3449 4886 3776
rect 4566 3213 4608 3449
rect 4844 3213 4886 3449
rect 4566 2752 4886 3213
rect 4566 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4814 2752
rect 4878 2688 4886 2752
rect 4566 2128 4886 2688
rect 5226 11042 5546 11472
rect 5226 10912 5268 11042
rect 5504 10912 5546 11042
rect 5226 10848 5234 10912
rect 5538 10848 5546 10912
rect 5226 10806 5268 10848
rect 5504 10806 5546 10848
rect 5226 9824 5546 10806
rect 5226 9760 5234 9824
rect 5298 9760 5314 9824
rect 5378 9760 5394 9824
rect 5458 9760 5474 9824
rect 5538 9760 5546 9824
rect 5226 8736 5546 9760
rect 5226 8672 5234 8736
rect 5298 8731 5314 8736
rect 5378 8731 5394 8736
rect 5458 8731 5474 8736
rect 5538 8672 5546 8736
rect 5226 8495 5268 8672
rect 5504 8495 5546 8672
rect 5226 7648 5546 8495
rect 5226 7584 5234 7648
rect 5298 7584 5314 7648
rect 5378 7584 5394 7648
rect 5458 7584 5474 7648
rect 5538 7584 5546 7648
rect 5226 6560 5546 7584
rect 5226 6496 5234 6560
rect 5298 6496 5314 6560
rect 5378 6496 5394 6560
rect 5458 6496 5474 6560
rect 5538 6496 5546 6560
rect 5226 6420 5546 6496
rect 5226 6184 5268 6420
rect 5504 6184 5546 6420
rect 5226 5472 5546 6184
rect 5226 5408 5234 5472
rect 5298 5408 5314 5472
rect 5378 5408 5394 5472
rect 5458 5408 5474 5472
rect 5538 5408 5546 5472
rect 5226 4384 5546 5408
rect 5226 4320 5234 4384
rect 5298 4320 5314 4384
rect 5378 4320 5394 4384
rect 5458 4320 5474 4384
rect 5538 4320 5546 4384
rect 5226 4109 5546 4320
rect 5226 3873 5268 4109
rect 5504 3873 5546 4109
rect 5226 3296 5546 3873
rect 5226 3232 5234 3296
rect 5298 3232 5314 3296
rect 5378 3232 5394 3296
rect 5458 3232 5474 3296
rect 5538 3232 5546 3296
rect 5226 2208 5546 3232
rect 5226 2144 5234 2208
rect 5298 2144 5314 2208
rect 5378 2144 5394 2208
rect 5458 2144 5474 2208
rect 5538 2144 5546 2208
rect 5226 2128 5546 2144
rect 6981 11456 7301 11472
rect 6981 11392 6989 11456
rect 7053 11392 7069 11456
rect 7133 11392 7149 11456
rect 7213 11392 7229 11456
rect 7293 11392 7301 11456
rect 6981 10382 7301 11392
rect 6981 10368 7023 10382
rect 7259 10368 7301 10382
rect 6981 10304 6989 10368
rect 7293 10304 7301 10368
rect 6981 10146 7023 10304
rect 7259 10146 7301 10304
rect 6981 9280 7301 10146
rect 6981 9216 6989 9280
rect 7053 9216 7069 9280
rect 7133 9216 7149 9280
rect 7213 9216 7229 9280
rect 7293 9216 7301 9280
rect 6981 8192 7301 9216
rect 6981 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7229 8192
rect 7293 8128 7301 8192
rect 6981 8071 7301 8128
rect 6981 7835 7023 8071
rect 7259 7835 7301 8071
rect 6981 7104 7301 7835
rect 6981 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7229 7104
rect 7293 7040 7301 7104
rect 6981 6016 7301 7040
rect 6981 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7229 6016
rect 7293 5952 7301 6016
rect 6981 5760 7301 5952
rect 6981 5524 7023 5760
rect 7259 5524 7301 5760
rect 6981 4928 7301 5524
rect 6981 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7229 4928
rect 7293 4864 7301 4928
rect 6981 3840 7301 4864
rect 6981 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7229 3840
rect 7293 3776 7301 3840
rect 6981 3449 7301 3776
rect 6981 3213 7023 3449
rect 7259 3213 7301 3449
rect 6981 2752 7301 3213
rect 6981 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7229 2752
rect 7293 2688 7301 2752
rect 6981 2128 7301 2688
rect 7641 11042 7961 11472
rect 7641 10912 7683 11042
rect 7919 10912 7961 11042
rect 7641 10848 7649 10912
rect 7953 10848 7961 10912
rect 7641 10806 7683 10848
rect 7919 10806 7961 10848
rect 7641 9824 7961 10806
rect 7641 9760 7649 9824
rect 7713 9760 7729 9824
rect 7793 9760 7809 9824
rect 7873 9760 7889 9824
rect 7953 9760 7961 9824
rect 7641 8736 7961 9760
rect 7641 8672 7649 8736
rect 7713 8731 7729 8736
rect 7793 8731 7809 8736
rect 7873 8731 7889 8736
rect 7953 8672 7961 8736
rect 7641 8495 7683 8672
rect 7919 8495 7961 8672
rect 7641 7648 7961 8495
rect 7641 7584 7649 7648
rect 7713 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7889 7648
rect 7953 7584 7961 7648
rect 7641 6560 7961 7584
rect 7641 6496 7649 6560
rect 7713 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7889 6560
rect 7953 6496 7961 6560
rect 7641 6420 7961 6496
rect 7641 6184 7683 6420
rect 7919 6184 7961 6420
rect 7641 5472 7961 6184
rect 7641 5408 7649 5472
rect 7713 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7889 5472
rect 7953 5408 7961 5472
rect 7641 4384 7961 5408
rect 7641 4320 7649 4384
rect 7713 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7889 4384
rect 7953 4320 7961 4384
rect 7641 4109 7961 4320
rect 7641 3873 7683 4109
rect 7919 3873 7961 4109
rect 7641 3296 7961 3873
rect 7641 3232 7649 3296
rect 7713 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7889 3296
rect 7953 3232 7961 3296
rect 7641 2208 7961 3232
rect 7641 2144 7649 2208
rect 7713 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7889 2208
rect 7953 2144 7961 2208
rect 7641 2128 7961 2144
rect 9396 11456 9716 11472
rect 9396 11392 9404 11456
rect 9468 11392 9484 11456
rect 9548 11392 9564 11456
rect 9628 11392 9644 11456
rect 9708 11392 9716 11456
rect 9396 10382 9716 11392
rect 9396 10368 9438 10382
rect 9674 10368 9716 10382
rect 9396 10304 9404 10368
rect 9708 10304 9716 10368
rect 9396 10146 9438 10304
rect 9674 10146 9716 10304
rect 9396 9280 9716 10146
rect 9396 9216 9404 9280
rect 9468 9216 9484 9280
rect 9548 9216 9564 9280
rect 9628 9216 9644 9280
rect 9708 9216 9716 9280
rect 9396 8192 9716 9216
rect 9396 8128 9404 8192
rect 9468 8128 9484 8192
rect 9548 8128 9564 8192
rect 9628 8128 9644 8192
rect 9708 8128 9716 8192
rect 9396 8071 9716 8128
rect 9396 7835 9438 8071
rect 9674 7835 9716 8071
rect 9396 7104 9716 7835
rect 9396 7040 9404 7104
rect 9468 7040 9484 7104
rect 9548 7040 9564 7104
rect 9628 7040 9644 7104
rect 9708 7040 9716 7104
rect 9396 6016 9716 7040
rect 9396 5952 9404 6016
rect 9468 5952 9484 6016
rect 9548 5952 9564 6016
rect 9628 5952 9644 6016
rect 9708 5952 9716 6016
rect 9396 5760 9716 5952
rect 9396 5524 9438 5760
rect 9674 5524 9716 5760
rect 9396 4928 9716 5524
rect 9396 4864 9404 4928
rect 9468 4864 9484 4928
rect 9548 4864 9564 4928
rect 9628 4864 9644 4928
rect 9708 4864 9716 4928
rect 9396 3840 9716 4864
rect 9396 3776 9404 3840
rect 9468 3776 9484 3840
rect 9548 3776 9564 3840
rect 9628 3776 9644 3840
rect 9708 3776 9716 3840
rect 9396 3449 9716 3776
rect 9396 3213 9438 3449
rect 9674 3213 9716 3449
rect 9396 2752 9716 3213
rect 9396 2688 9404 2752
rect 9468 2688 9484 2752
rect 9548 2688 9564 2752
rect 9628 2688 9644 2752
rect 9708 2688 9716 2752
rect 9396 2128 9716 2688
rect 10056 11042 10376 11472
rect 10056 10912 10098 11042
rect 10334 10912 10376 11042
rect 10056 10848 10064 10912
rect 10368 10848 10376 10912
rect 10056 10806 10098 10848
rect 10334 10806 10376 10848
rect 10056 9824 10376 10806
rect 10056 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10376 9824
rect 10056 8736 10376 9760
rect 10056 8672 10064 8736
rect 10128 8731 10144 8736
rect 10208 8731 10224 8736
rect 10288 8731 10304 8736
rect 10368 8672 10376 8736
rect 10056 8495 10098 8672
rect 10334 8495 10376 8672
rect 10056 7648 10376 8495
rect 10056 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10376 7648
rect 10056 6560 10376 7584
rect 10056 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10376 6560
rect 10056 6420 10376 6496
rect 10056 6184 10098 6420
rect 10334 6184 10376 6420
rect 10056 5472 10376 6184
rect 10056 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10376 5472
rect 10056 4384 10376 5408
rect 10056 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10376 4384
rect 10056 4109 10376 4320
rect 10056 3873 10098 4109
rect 10334 3873 10376 4109
rect 10056 3296 10376 3873
rect 10056 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10376 3296
rect 10056 2208 10376 3232
rect 10056 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10376 2208
rect 10056 2128 10376 2144
<< via4 >>
rect 2193 10368 2429 10382
rect 2193 10304 2223 10368
rect 2223 10304 2239 10368
rect 2239 10304 2303 10368
rect 2303 10304 2319 10368
rect 2319 10304 2383 10368
rect 2383 10304 2399 10368
rect 2399 10304 2429 10368
rect 2193 10146 2429 10304
rect 2193 7835 2429 8071
rect 2193 5524 2429 5760
rect 2193 3213 2429 3449
rect 2853 10912 3089 11042
rect 2853 10848 2883 10912
rect 2883 10848 2899 10912
rect 2899 10848 2963 10912
rect 2963 10848 2979 10912
rect 2979 10848 3043 10912
rect 3043 10848 3059 10912
rect 3059 10848 3089 10912
rect 2853 10806 3089 10848
rect 2853 8672 2883 8731
rect 2883 8672 2899 8731
rect 2899 8672 2963 8731
rect 2963 8672 2979 8731
rect 2979 8672 3043 8731
rect 3043 8672 3059 8731
rect 3059 8672 3089 8731
rect 2853 8495 3089 8672
rect 2853 6184 3089 6420
rect 2853 3873 3089 4109
rect 4608 10368 4844 10382
rect 4608 10304 4638 10368
rect 4638 10304 4654 10368
rect 4654 10304 4718 10368
rect 4718 10304 4734 10368
rect 4734 10304 4798 10368
rect 4798 10304 4814 10368
rect 4814 10304 4844 10368
rect 4608 10146 4844 10304
rect 4608 7835 4844 8071
rect 4608 5524 4844 5760
rect 4608 3213 4844 3449
rect 5268 10912 5504 11042
rect 5268 10848 5298 10912
rect 5298 10848 5314 10912
rect 5314 10848 5378 10912
rect 5378 10848 5394 10912
rect 5394 10848 5458 10912
rect 5458 10848 5474 10912
rect 5474 10848 5504 10912
rect 5268 10806 5504 10848
rect 5268 8672 5298 8731
rect 5298 8672 5314 8731
rect 5314 8672 5378 8731
rect 5378 8672 5394 8731
rect 5394 8672 5458 8731
rect 5458 8672 5474 8731
rect 5474 8672 5504 8731
rect 5268 8495 5504 8672
rect 5268 6184 5504 6420
rect 5268 3873 5504 4109
rect 7023 10368 7259 10382
rect 7023 10304 7053 10368
rect 7053 10304 7069 10368
rect 7069 10304 7133 10368
rect 7133 10304 7149 10368
rect 7149 10304 7213 10368
rect 7213 10304 7229 10368
rect 7229 10304 7259 10368
rect 7023 10146 7259 10304
rect 7023 7835 7259 8071
rect 7023 5524 7259 5760
rect 7023 3213 7259 3449
rect 7683 10912 7919 11042
rect 7683 10848 7713 10912
rect 7713 10848 7729 10912
rect 7729 10848 7793 10912
rect 7793 10848 7809 10912
rect 7809 10848 7873 10912
rect 7873 10848 7889 10912
rect 7889 10848 7919 10912
rect 7683 10806 7919 10848
rect 7683 8672 7713 8731
rect 7713 8672 7729 8731
rect 7729 8672 7793 8731
rect 7793 8672 7809 8731
rect 7809 8672 7873 8731
rect 7873 8672 7889 8731
rect 7889 8672 7919 8731
rect 7683 8495 7919 8672
rect 7683 6184 7919 6420
rect 7683 3873 7919 4109
rect 9438 10368 9674 10382
rect 9438 10304 9468 10368
rect 9468 10304 9484 10368
rect 9484 10304 9548 10368
rect 9548 10304 9564 10368
rect 9564 10304 9628 10368
rect 9628 10304 9644 10368
rect 9644 10304 9674 10368
rect 9438 10146 9674 10304
rect 9438 7835 9674 8071
rect 9438 5524 9674 5760
rect 9438 3213 9674 3449
rect 10098 10912 10334 11042
rect 10098 10848 10128 10912
rect 10128 10848 10144 10912
rect 10144 10848 10208 10912
rect 10208 10848 10224 10912
rect 10224 10848 10288 10912
rect 10288 10848 10304 10912
rect 10304 10848 10334 10912
rect 10098 10806 10334 10848
rect 10098 8672 10128 8731
rect 10128 8672 10144 8731
rect 10144 8672 10208 8731
rect 10208 8672 10224 8731
rect 10224 8672 10288 8731
rect 10288 8672 10304 8731
rect 10304 8672 10334 8731
rect 10098 8495 10334 8672
rect 10098 6184 10334 6420
rect 10098 3873 10334 4109
<< metal5 >>
rect 1056 11042 10812 11084
rect 1056 10806 2853 11042
rect 3089 10806 5268 11042
rect 5504 10806 7683 11042
rect 7919 10806 10098 11042
rect 10334 10806 10812 11042
rect 1056 10764 10812 10806
rect 1056 10382 10812 10424
rect 1056 10146 2193 10382
rect 2429 10146 4608 10382
rect 4844 10146 7023 10382
rect 7259 10146 9438 10382
rect 9674 10146 10812 10382
rect 1056 10104 10812 10146
rect 1056 8731 10812 8773
rect 1056 8495 2853 8731
rect 3089 8495 5268 8731
rect 5504 8495 7683 8731
rect 7919 8495 10098 8731
rect 10334 8495 10812 8731
rect 1056 8453 10812 8495
rect 1056 8071 10812 8113
rect 1056 7835 2193 8071
rect 2429 7835 4608 8071
rect 4844 7835 7023 8071
rect 7259 7835 9438 8071
rect 9674 7835 10812 8071
rect 1056 7793 10812 7835
rect 1056 6420 10812 6462
rect 1056 6184 2853 6420
rect 3089 6184 5268 6420
rect 5504 6184 7683 6420
rect 7919 6184 10098 6420
rect 10334 6184 10812 6420
rect 1056 6142 10812 6184
rect 1056 5760 10812 5802
rect 1056 5524 2193 5760
rect 2429 5524 4608 5760
rect 4844 5524 7023 5760
rect 7259 5524 9438 5760
rect 9674 5524 10812 5760
rect 1056 5482 10812 5524
rect 1056 4109 10812 4151
rect 1056 3873 2853 4109
rect 3089 3873 5268 4109
rect 5504 3873 7683 4109
rect 7919 3873 10098 4109
rect 10334 3873 10812 4109
rect 1056 3831 10812 3873
rect 1056 3449 10812 3491
rect 1056 3213 2193 3449
rect 2429 3213 4608 3449
rect 4844 3213 7023 3449
rect 7259 3213 9438 3449
rect 9674 3213 10812 3449
rect 1056 3171 10812 3213
use sky130_fd_sc_hd__or3b_1  _049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 4232 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 5152 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5980 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _053_
timestamp 1717180972
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1717180972
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1717180972
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 4416 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _058_
timestamp 1717180972
transform 1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _059_
timestamp 1717180972
transform 1 0 3772 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _060_
timestamp 1717180972
transform -1 0 3772 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _063_
timestamp 1717180972
transform -1 0 10396 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _065_
timestamp 1717180972
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10028 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 8096 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _071_
timestamp 1717180972
transform -1 0 8740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 7636 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1717180972
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _074_
timestamp 1717180972
transform 1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _075_
timestamp 1717180972
transform 1 0 8004 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _076_
timestamp 1717180972
transform 1 0 3128 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _077_
timestamp 1717180972
transform -1 0 4416 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _078_
timestamp 1717180972
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _079_
timestamp 1717180972
transform -1 0 3680 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _080_
timestamp 1717180972
transform -1 0 2208 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _082_
timestamp 1717180972
transform -1 0 2392 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _083_
timestamp 1717180972
transform -1 0 2484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1717180972
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9936 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _087_
timestamp 1717180972
transform 1 0 8372 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _088_
timestamp 1717180972
transform -1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _089_
timestamp 1717180972
transform -1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1717180972
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1717180972
transform -1 0 8740 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1717180972
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _093_
timestamp 1717180972
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _095_
timestamp 1717180972
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _096_
timestamp 1717180972
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7268 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 6072 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _099_
timestamp 1717180972
transform 1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _103_
timestamp 1717180972
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp 1717180972
transform 1 0 8464 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp 1717180972
transform 1 0 9016 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _107_
timestamp 1717180972
transform 1 0 7084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 1717180972
transform 1 0 7636 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _109_
timestamp 1717180972
transform 1 0 3772 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _110_
timestamp 1717180972
transform 1 0 1932 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _111_
timestamp 1717180972
transform -1 0 5796 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp 1717180972
transform 1 0 3772 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp 1717180972
transform 1 0 1564 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp 1717180972
transform 1 0 1656 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _115_
timestamp 1717180972
transform 1 0 9016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _116_
timestamp 1717180972
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 1717180972
transform 1 0 5244 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 1717180972
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp 1717180972
transform 1 0 5520 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _120_
timestamp 1717180972
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 1717180972
transform -1 0 5704 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 1717180972
transform 1 0 6256 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _123_
timestamp 1717180972
transform 1 0 9016 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 1717180972
transform 1 0 7912 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5336 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1717180972
transform -1 0 6256 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1717180972
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 1717180972
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1717180972
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1717180972
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_11
timestamp 1717180972
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_29
timestamp 1717180972
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1717180972
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1717180972
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1717180972
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1717180972
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_96
timestamp 1717180972
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1717180972
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1717180972
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1717180972
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1717180972
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 1717180972
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 1717180972
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_43
timestamp 1717180972
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1717180972
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1717180972
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1717180972
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1717180972
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_97
timestamp 1717180972
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_101
timestamp 1717180972
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1717180972
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1717180972
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1717180972
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1717180972
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_43
timestamp 1717180972
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_55
timestamp 1717180972
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1717180972
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1717180972
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_29
timestamp 1717180972
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1717180972
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1717180972
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_77
timestamp 1717180972
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_96
timestamp 1717180972
transform 1 0 9936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1717180972
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 1717180972
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_40
timestamp 1717180972
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_44
timestamp 1717180972
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_68
timestamp 1717180972
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_76
timestamp 1717180972
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1717180972
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1717180972
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_99
timestamp 1717180972
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1717180972
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1717180972
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 1717180972
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1717180972
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1717180972
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_61
timestamp 1717180972
transform 1 0 6716 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_69
timestamp 1717180972
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_75
timestamp 1717180972
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1717180972
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1717180972
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1717180972
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1717180972
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_32
timestamp 1717180972
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_66
timestamp 1717180972
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1717180972
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1717180972
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_26
timestamp 1717180972
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_49
timestamp 1717180972
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 1717180972
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_86
timestamp 1717180972
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_101
timestamp 1717180972
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1717180972
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_12
timestamp 1717180972
transform 1 0 2208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_20
timestamp 1717180972
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1717180972
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 1717180972
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1717180972
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1717180972
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_100
timestamp 1717180972
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1717180972
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_25
timestamp 1717180972
transform 1 0 3404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_29
timestamp 1717180972
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1717180972
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1717180972
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1717180972
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_62
timestamp 1717180972
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_71
timestamp 1717180972
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_90
timestamp 1717180972
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1717180972
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1717180972
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1717180972
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1717180972
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1717180972
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_42
timestamp 1717180972
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_52
timestamp 1717180972
transform 1 0 5888 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_58
timestamp 1717180972
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_70
timestamp 1717180972
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1717180972
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1717180972
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1717180972
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1717180972
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_44
timestamp 1717180972
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1717180972
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_72
timestamp 1717180972
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_82
timestamp 1717180972
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1717180972
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1717180972
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1717180972
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1717180972
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1717180972
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_96
timestamp 1717180972
transform 1 0 9936 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_6
timestamp 1717180972
transform 1 0 1656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_12
timestamp 1717180972
transform 1 0 2208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_28
timestamp 1717180972
transform 1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1717180972
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_71
timestamp 1717180972
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_87
timestamp 1717180972
transform 1 0 9108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1717180972
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_15
timestamp 1717180972
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1717180972
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_29
timestamp 1717180972
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_40
timestamp 1717180972
transform 1 0 4784 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_52
timestamp 1717180972
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_57
timestamp 1717180972
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_68
timestamp 1717180972
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1717180972
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1717180972
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_92
timestamp 1717180972
transform 1 0 9568 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_100
timestamp 1717180972
transform 1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1717180972
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1717180972
transform -1 0 8740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1717180972
transform 1 0 7268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1717180972
transform -1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1717180972
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1717180972
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1717180972
transform -1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1717180972
transform -1 0 4784 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1717180972
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1717180972
transform -1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1717180972
transform -1 0 9936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1717180972
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1717180972
transform -1 0 3128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1717180972
transform -1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold17
timestamp 1717180972
transform -1 0 5336 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1717180972
transform 1 0 4048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  hold20
timestamp 1717180972
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1717180972
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold22
timestamp 1717180972
transform 1 0 4140 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1717180972
transform 1 0 5152 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1717180972
transform -1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold25
timestamp 1717180972
transform -1 0 4140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1717180972
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1717180972
transform -1 0 10396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1717180972
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1717180972
transform -1 0 8648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1717180972
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1717180972
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1717180972
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1717180972
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1717180972
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1717180972
transform 1 0 9016 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1717180972
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1717180972
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1717180972
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1717180972
transform -1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1717180972
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1717180972
transform -1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1717180972
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1717180972
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1717180972
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1717180972
transform -1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1717180972
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1717180972
transform -1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1717180972
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1717180972
transform -1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1717180972
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1717180972
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1717180972
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1717180972
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1717180972
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1717180972
transform -1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1717180972
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1717180972
transform -1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1717180972
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1717180972
transform -1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1717180972
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1717180972
transform -1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1717180972
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1717180972
transform -1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1717180972
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1717180972
transform -1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1717180972
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1717180972
transform -1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1717180972
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1717180972
transform -1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1717180972
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1717180972
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1717180972
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1717180972
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1717180972
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1717180972
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1717180972
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1717180972
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1717180972
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1717180972
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1717180972
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1717180972
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1717180972
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1717180972
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1717180972
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1717180972
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1717180972
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1717180972
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1717180972
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1717180972
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1717180972
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1717180972
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1717180972
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1717180972
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1717180972
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1717180972
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1717180972
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 2811 2128 3131 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5226 2128 5546 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7641 2128 7961 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10056 2128 10376 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3831 10812 4151 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6142 10812 6462 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8453 10812 8773 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10764 10812 11084 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2151 2128 2471 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4566 2128 4886 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6981 2128 7301 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9396 2128 9716 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3171 10812 3491 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5482 10812 5802 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7793 10812 8113 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 10104 10812 10424 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 11154 3272 11954 3392 0 FreeSans 480 0 0 0 percentage[0]
port 3 nsew signal input
flabel metal3 s 11154 10344 11954 10464 0 FreeSans 480 0 0 0 percentage[1]
port 4 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 s_in_lines[0]
port 5 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 s_in_lines[1]
port 6 nsew signal input
flabel metal2 s 2962 13298 3018 14098 0 FreeSans 224 90 0 0 s_out_lines[0]
port 7 nsew signal tristate
flabel metal2 s 8942 13298 8998 14098 0 FreeSans 224 90 0 0 s_out_lines[1]
port 8 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 start
port 9 nsew signal input
rlabel metal1 5934 10880 5934 10880 0 VGND
rlabel metal1 5934 11424 5934 11424 0 VPWR
rlabel metal1 7682 7514 7682 7514 0 CTRLPTH1.done
rlabel metal1 6578 8568 6578 8568 0 CTRLPTH1.state\[0\]
rlabel metal1 5428 8942 5428 8942 0 CTRLPTH1.state\[1\]
rlabel metal1 7360 10574 7360 10574 0 CTRLPTH1.state\[2\]
rlabel metal1 10626 9010 10626 9010 0 DTPTH1.PS1.count\[0\]
rlabel metal2 9338 8058 9338 8058 0 DTPTH1.PS1.count\[1\]
rlabel metal1 3496 6766 3496 6766 0 DTPTH1.RS1.RNG1.TFF1.Q
rlabel metal1 4048 8466 4048 8466 0 DTPTH1.RS1.RNG1.TFF2.Q
rlabel metal1 5428 6834 5428 6834 0 DTPTH1.RS1.RNG1.TFF3.Q
rlabel metal2 4002 5508 4002 5508 0 DTPTH1.RS1.RNG1.TFF4.Q
rlabel metal1 3956 4658 3956 4658 0 DTPTH1.RS1.RNG1.TFF5.Q
rlabel metal1 5612 2618 5612 2618 0 DTPTH1.RS1.RNG1.TFF6.Q
rlabel metal1 4370 3468 4370 3468 0 DTPTH1.RS1.RNG1.TFF7.Q
rlabel metal1 4738 6154 4738 6154 0 DTPTH1.RS1.RNG1.b0
rlabel metal1 6210 5270 6210 5270 0 DTPTH1.RS1.RNG1.b1
rlabel metal1 5106 4046 5106 4046 0 DTPTH1.RS1.RNG1.b2
rlabel metal1 7958 4046 7958 4046 0 DTPTH1.RS1.RNG1.r_num\[0\]
rlabel metal1 8786 3434 8786 3434 0 DTPTH1.RS1.RNG1.r_num\[1\]
rlabel metal1 7866 5882 7866 5882 0 DTPTH1.RS1.RNG1.r_num\[2\]
rlabel metal1 10304 7446 10304 7446 0 DTPTH1.RS1.counter\[0\]
rlabel metal1 9522 6868 9522 6868 0 DTPTH1.RS1.counter\[1\]
rlabel metal1 10120 4658 10120 4658 0 DTPTH1.RS1.s_comb\[0\]
rlabel metal1 10212 3706 10212 3706 0 DTPTH1.RS1.s_comb\[1\]
rlabel metal2 8602 4148 8602 4148 0 DTPTH1.RS1.s_comb\[2\]
rlabel metal1 9292 2482 9292 2482 0 DTPTH1.RS1.s_comb\[3\]
rlabel metal1 5435 7378 5435 7378 0 _000_
rlabel metal1 4646 9486 4646 9486 0 _001_
rlabel metal2 3174 4352 3174 4352 0 _002_
rlabel metal1 6568 7378 6568 7378 0 _003_
rlabel metal1 9752 4794 9752 4794 0 _004_
rlabel metal1 9246 3060 9246 3060 0 _005_
rlabel metal1 7268 4250 7268 4250 0 _006_
rlabel metal1 8004 2618 8004 2618 0 _007_
rlabel metal1 4048 2346 4048 2346 0 _008_
rlabel metal1 2484 5134 2484 5134 0 _009_
rlabel metal1 3864 5746 3864 5746 0 _010_
rlabel metal1 2507 6766 2507 6766 0 _011_
rlabel metal1 1748 8058 1748 8058 0 _012_
rlabel metal2 1978 7140 1978 7140 0 _013_
rlabel metal1 8970 6392 8970 6392 0 _014_
rlabel metal1 7636 6426 7636 6426 0 _015_
rlabel metal1 3894 9962 3894 9962 0 _016_
rlabel metal1 5581 10710 5581 10710 0 _017_
rlabel metal2 6578 9826 6578 9826 0 _018_
rlabel metal1 9425 9622 9425 9622 0 _019_
rlabel via1 8229 8466 8229 8466 0 _020_
rlabel metal1 6944 9554 6944 9554 0 _021_
rlabel metal1 3956 9010 3956 9010 0 _022_
rlabel metal1 7130 10642 7130 10642 0 _023_
rlabel metal1 9890 10064 9890 10064 0 _024_
rlabel metal1 8372 9554 8372 9554 0 _025_
rlabel metal2 7406 10302 7406 10302 0 _026_
rlabel metal1 7866 8840 7866 8840 0 _027_
rlabel metal1 10258 7174 10258 7174 0 _028_
rlabel metal1 7544 7174 7544 7174 0 _029_
rlabel metal1 6118 7378 6118 7378 0 _030_
rlabel metal1 9062 4250 9062 4250 0 _031_
rlabel metal1 8970 8874 8970 8874 0 _032_
rlabel metal1 8326 2448 8326 2448 0 _033_
rlabel metal1 8372 2550 8372 2550 0 _034_
rlabel metal1 8464 3638 8464 3638 0 _035_
rlabel metal1 2346 5746 2346 5746 0 _036_
rlabel metal2 1886 6358 1886 6358 0 _037_
rlabel metal1 8142 7344 8142 7344 0 _038_
rlabel metal1 9384 7514 9384 7514 0 _039_
rlabel metal1 10074 6834 10074 6834 0 _040_
rlabel metal1 10166 5712 10166 5712 0 _041_
rlabel metal1 9936 5542 9936 5542 0 _042_
rlabel metal2 8326 7616 8326 7616 0 _043_
rlabel metal1 8648 7514 8648 7514 0 _044_
rlabel metal1 5750 10608 5750 10608 0 _045_
rlabel metal1 3542 10234 3542 10234 0 _046_
rlabel metal2 8418 10472 8418 10472 0 _047_
rlabel metal2 8142 10472 8142 10472 0 _048_
rlabel metal3 1671 3332 1671 3332 0 clk
rlabel metal1 6440 6630 6440 6630 0 clknet_0_clk
rlabel metal1 1794 3570 1794 3570 0 clknet_1_0__leaf_clk
rlabel metal2 1610 7922 1610 7922 0 clknet_1_1__leaf_clk
rlabel metal1 10074 10234 10074 10234 0 net1
rlabel metal2 7498 4352 7498 4352 0 net10
rlabel metal1 7493 3434 7493 3434 0 net11
rlabel metal1 8740 2414 8740 2414 0 net12
rlabel metal1 5704 9146 5704 9146 0 net13
rlabel metal2 6026 9146 6026 9146 0 net14
rlabel metal1 4455 2346 4455 2346 0 net15
rlabel metal1 4462 9554 4462 9554 0 net16
rlabel metal2 3358 10608 3358 10608 0 net17
rlabel metal1 5014 9146 5014 9146 0 net18
rlabel metal1 9614 4590 9614 4590 0 net19
rlabel metal1 9200 10030 9200 10030 0 net2
rlabel metal1 9011 5270 9011 5270 0 net20
rlabel metal1 3680 3026 3680 3026 0 net21
rlabel metal1 2162 3162 2162 3162 0 net22
rlabel metal1 7360 9486 7360 9486 0 net23
rlabel metal2 3358 6511 3358 6511 0 net24
rlabel metal1 5474 5304 5474 5304 0 net25
rlabel metal1 5106 5542 5106 5542 0 net26
rlabel metal1 1886 7854 1886 7854 0 net27
rlabel metal2 5842 5916 5842 5916 0 net28
rlabel metal1 3818 4114 3818 4114 0 net29
rlabel metal1 3174 2618 3174 2618 0 net3
rlabel metal1 5651 3706 5651 3706 0 net30
rlabel metal1 3956 3706 3956 3706 0 net31
rlabel metal1 3726 7922 3726 7922 0 net32
rlabel metal1 9752 8942 9752 8942 0 net33
rlabel metal1 8694 6256 8694 6256 0 net34
rlabel metal1 8786 6970 8786 6970 0 net35
rlabel metal1 8004 6290 8004 6290 0 net36
rlabel metal1 8326 2278 8326 2278 0 net4
rlabel metal1 1610 10132 1610 10132 0 net5
rlabel metal2 3174 10914 3174 10914 0 net6
rlabel metal1 9108 10778 9108 10778 0 net7
rlabel metal1 8464 2822 8464 2822 0 net8
rlabel metal2 9890 3298 9890 3298 0 net9
rlabel metal1 10672 3026 10672 3026 0 percentage[0]
rlabel metal1 10672 10642 10672 10642 0 percentage[1]
rlabel metal2 2990 823 2990 823 0 s_in_lines[0]
rlabel metal2 8970 1027 8970 1027 0 s_in_lines[1]
rlabel metal1 3128 11322 3128 11322 0 s_out_lines[0]
rlabel metal1 9108 11322 9108 11322 0 s_out_lines[1]
rlabel metal3 820 10404 820 10404 0 start
<< properties >>
string FIXED_BBOX 0 0 11954 14098
<< end >>
