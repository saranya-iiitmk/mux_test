magic
tech sky130A
magscale 1 2
timestamp 1717180972
<< dnwell >>
rect 5296 -6592 8535 -5514
<< nwell >>
rect 5847 -2455 6881 -2287
rect 5848 -2814 6872 -2455
rect 5848 -2818 6536 -2814
rect 5848 -2852 6551 -2818
rect 6594 -2852 6872 -2814
rect 5848 -2970 6872 -2852
rect 5216 -5720 8620 -5434
rect 5216 -6386 5502 -5720
rect 8318 -6386 8620 -5720
rect 5216 -6672 8620 -6386
<< pwell >>
rect 6762 -6202 6828 -6192
rect 7168 -6200 7234 -6190
rect 6148 -6344 6250 -6310
rect 6548 -6344 6650 -6310
rect 6938 -6342 7040 -6308
rect 7340 -6342 7442 -6308
rect 7748 -6342 7850 -6308
<< psubdiff >>
rect 6148 -6344 6250 -6310
rect 6548 -6344 6650 -6310
rect 6938 -6342 7040 -6308
rect 7340 -6342 7442 -6308
rect 7748 -6342 7850 -6308
<< nsubdiff >>
rect 5253 -5491 8567 -5471
rect 5253 -5525 5333 -5491
rect 8487 -5525 8567 -5491
rect 5253 -5545 8567 -5525
rect 5253 -5551 5327 -5545
rect 5253 -6555 5273 -5551
rect 5307 -6555 5327 -5551
rect 8493 -5551 8567 -5545
rect 5253 -6561 5327 -6555
rect 8493 -6555 8513 -5551
rect 8547 -6555 8567 -5551
rect 8493 -6561 8567 -6555
rect 5253 -6581 8567 -6561
rect 5253 -6615 5333 -6581
rect 8487 -6615 8567 -6581
rect 5253 -6635 8567 -6615
<< nsubdiffcont >>
rect 5333 -5525 8487 -5491
rect 5273 -6555 5307 -5551
rect 8513 -6555 8547 -5551
rect 5333 -6615 8487 -6581
<< poly >>
rect 5888 -2391 5963 -2374
rect 5888 -2426 5909 -2391
rect 5943 -2396 5963 -2391
rect 6492 -2387 6559 -2370
rect 5943 -2426 6235 -2396
rect 5888 -2443 5963 -2426
rect 6204 -2484 6235 -2426
rect 6492 -2422 6510 -2387
rect 6544 -2422 6559 -2387
rect 6492 -2439 6559 -2422
rect 6204 -2514 6322 -2484
rect 6204 -2584 6234 -2514
rect 6292 -2580 6322 -2514
rect 6506 -2594 6536 -2439
rect 6594 -2919 6624 -2814
rect 6576 -2929 6642 -2919
rect 6576 -2963 6592 -2929
rect 6626 -2963 6642 -2929
rect 6576 -2973 6642 -2963
rect 4943 -5612 5020 -5599
rect 4943 -5647 4965 -5612
rect 5000 -5647 5020 -5612
rect 4943 -5663 5020 -5647
rect 4943 -5700 4973 -5663
rect 6762 -6202 6828 -6192
rect 7168 -6200 7234 -6190
<< polycont >>
rect 5909 -2426 5943 -2391
rect 6510 -2422 6544 -2387
rect 6592 -2963 6626 -2929
rect 4965 -5647 5000 -5612
<< locali >>
rect 5888 -2389 5963 -2374
rect 5888 -2426 5909 -2389
rect 5944 -2426 5963 -2389
rect 5888 -2443 5963 -2426
rect 6492 -2387 6559 -2370
rect 6492 -2422 6510 -2387
rect 6544 -2422 6559 -2387
rect 6492 -2439 6559 -2422
rect 6026 -2556 6582 -2522
rect 6026 -5173 6060 -2556
rect 6246 -2590 6280 -2556
rect 6548 -2590 6582 -2556
rect 6592 -2929 6626 -2913
rect 6592 -2979 6626 -2963
rect 4985 -5207 6060 -5173
rect 4985 -5599 5019 -5207
rect 5273 -5525 5333 -5491
rect 8487 -5525 8547 -5491
rect 5273 -5551 5307 -5525
rect 4943 -5612 5020 -5599
rect 4943 -5647 4965 -5612
rect 5000 -5647 5020 -5612
rect 4943 -5663 5020 -5647
rect 4985 -5720 5019 -5663
rect 4796 -5833 4899 -5825
rect 4796 -5860 4903 -5833
rect 8513 -5551 8547 -5525
rect 5808 -5705 5842 -5694
rect 5808 -5796 5842 -5739
rect 6004 -6092 6362 -6036
rect 7628 -6096 7986 -6040
rect 6148 -6344 6250 -6310
rect 6548 -6344 6650 -6310
rect 6938 -6342 7040 -6308
rect 7340 -6342 7442 -6308
rect 7748 -6342 7850 -6308
rect 5273 -6581 5307 -6555
rect 8513 -6581 8547 -6555
rect 5273 -6615 5333 -6581
rect 8487 -6615 8547 -6581
<< viali >>
rect 5909 -2391 5944 -2389
rect 5909 -2426 5943 -2391
rect 5943 -2426 5944 -2391
rect 6510 -2422 6544 -2387
rect 6592 -2963 6626 -2929
rect 5808 -5739 5842 -5705
<< metal1 >>
rect 5888 -2389 5963 -2374
rect 6492 -2386 6559 -2370
rect 5888 -2426 5909 -2389
rect 5944 -2426 5963 -2389
rect 5888 -2443 5963 -2426
rect 6328 -2387 6559 -2386
rect 6328 -2422 6510 -2387
rect 6544 -2422 6559 -2387
rect 6328 -2426 6559 -2422
rect 5905 -2880 5943 -2443
rect 6328 -2594 6374 -2426
rect 6492 -2439 6559 -2426
rect 6158 -2880 6192 -2747
rect 5905 -2913 6194 -2880
rect 6158 -5138 6192 -2913
rect 6334 -3442 6368 -2755
rect 6640 -2769 6860 -2735
rect 6460 -2929 6494 -2770
rect 6586 -2929 6632 -2917
rect 6460 -2963 6592 -2929
rect 6626 -2963 6632 -2929
rect 6460 -3100 6494 -2963
rect 6586 -2975 6632 -2963
rect 6451 -3106 6503 -3100
rect 6451 -3164 6503 -3158
rect 6286 -3454 6376 -3442
rect 6286 -3514 6292 -3454
rect 6358 -3514 6376 -3454
rect 6286 -3526 6376 -3514
rect 6334 -4880 6368 -3526
rect 6826 -4183 6860 -2769
rect 7433 -4183 7654 -4156
rect 6825 -4188 7654 -4183
rect 6825 -4311 7475 -4188
rect 6584 -4375 6636 -4369
rect 6584 -4433 6636 -4427
rect 6334 -4886 6390 -4880
rect 6334 -4948 6390 -4942
rect 6149 -5144 6201 -5138
rect 6149 -5202 6201 -5196
rect 5808 -5699 5842 -5351
rect 6593 -5644 6627 -4433
rect 6826 -5240 6860 -4311
rect 7433 -4339 7475 -4311
rect 7618 -4339 7654 -4188
rect 7433 -4378 7654 -4339
rect 6826 -5274 8267 -5240
rect 6593 -5678 8025 -5644
rect 5796 -5705 5854 -5699
rect 5796 -5739 5808 -5705
rect 5842 -5739 5854 -5705
rect 5796 -5745 5854 -5739
rect 6483 -5853 7025 -5799
rect 4897 -6097 4931 -5883
rect 5950 -5942 6016 -5882
rect 6356 -5942 6422 -5882
rect 6490 -6056 6530 -5853
rect 6630 -5968 6636 -5916
rect 6688 -5968 6694 -5916
rect 6762 -5942 6826 -5884
rect 5610 -6109 5958 -6076
rect 6418 -6096 6530 -6056
rect 6639 -6042 6685 -5968
rect 6971 -6042 7025 -5853
rect 7170 -5938 7234 -5880
rect 7266 -5894 7322 -5888
rect 7266 -6030 7322 -5950
rect 6639 -6088 6766 -6042
rect 6822 -6096 7176 -6042
rect 7228 -6086 7322 -6030
rect 7506 -6044 7540 -5678
rect 7991 -5884 8025 -5678
rect 7574 -5940 7638 -5886
rect 7978 -5940 8042 -5884
rect 8233 -5997 8267 -5274
rect 8049 -6031 8267 -5997
rect 7506 -6078 7578 -6044
rect 5610 -7000 5643 -6109
rect 5925 -6198 5958 -6109
rect 5925 -6209 6016 -6198
rect 6356 -6209 6422 -6198
rect 5925 -6242 6422 -6209
rect 5950 -6258 6016 -6242
rect 6356 -6258 6422 -6242
rect 6756 -6200 6834 -6198
rect 6756 -6256 6762 -6200
rect 6828 -6256 6834 -6200
rect 6377 -6319 6410 -6258
rect 6756 -6262 6834 -6256
rect 7166 -6200 7234 -6198
rect 7166 -6252 7174 -6200
rect 7226 -6252 7234 -6200
rect 7574 -6252 7638 -6196
rect 7166 -6258 7234 -6252
rect 7593 -6319 7626 -6252
rect 7980 -6254 8040 -6198
rect 6377 -6352 7626 -6319
rect 5890 -6769 5924 -6722
rect 6288 -6769 6294 -6760
rect 5890 -6803 6294 -6769
rect 5890 -6804 5924 -6803
rect 6288 -6812 6294 -6803
rect 6346 -6812 6352 -6760
rect 7146 -6880 7227 -6872
rect 7146 -6892 7158 -6880
rect 6468 -6934 7158 -6892
rect 7216 -6934 7227 -6880
rect 6468 -6946 7227 -6934
rect 4895 -7036 5643 -7000
rect 4895 -7037 5642 -7036
<< via1 >>
rect 6451 -3158 6503 -3106
rect 6292 -3514 6358 -3454
rect 6584 -4427 6636 -4375
rect 6334 -4942 6390 -4886
rect 6149 -5196 6201 -5144
rect 7475 -4339 7618 -4188
rect 6636 -5968 6688 -5916
rect 7266 -5950 7322 -5894
rect 6762 -6256 6828 -6200
rect 7174 -6252 7226 -6200
rect 6294 -6812 6346 -6760
rect 7158 -6934 7216 -6880
<< metal2 >>
rect 6436 -3102 6520 -3090
rect 6436 -3162 6447 -3102
rect 6507 -3162 6520 -3102
rect 6436 -3174 6520 -3162
rect 6286 -3454 6376 -3442
rect 6286 -3514 6292 -3454
rect 6358 -3514 6376 -3454
rect 6286 -3526 6376 -3514
rect 7433 -4188 7654 -4156
rect 7433 -4339 7475 -4188
rect 7618 -4339 7654 -4188
rect 6568 -4371 6651 -4356
rect 6568 -4431 6580 -4371
rect 6640 -4431 6651 -4371
rect 7433 -4378 7654 -4339
rect 6568 -4448 6651 -4431
rect 6328 -4942 6334 -4886
rect 6390 -4942 7322 -4886
rect 6151 -5144 6197 -5141
rect 6143 -5196 6149 -5144
rect 6201 -5157 6207 -5144
rect 6201 -5196 6545 -5157
rect 6151 -5203 6545 -5196
rect 6151 -5204 6197 -5203
rect 6499 -5749 6545 -5203
rect 6499 -5795 6685 -5749
rect 6639 -5910 6685 -5795
rect 7266 -5894 7322 -4942
rect 6636 -5916 6688 -5910
rect 7260 -5950 7266 -5894
rect 7322 -5950 7328 -5894
rect 6636 -5974 6688 -5968
rect 6756 -6200 6834 -6198
rect 6756 -6256 6762 -6200
rect 6828 -6256 6834 -6200
rect 7168 -6252 7174 -6200
rect 7226 -6252 7234 -6200
rect 7168 -6256 7234 -6252
rect 6756 -6262 6834 -6256
rect 6770 -6286 6814 -6262
rect 6294 -6760 6346 -6754
rect 6775 -6773 6805 -6286
rect 6346 -6803 6805 -6773
rect 6294 -6818 6346 -6812
rect 7186 -6872 7218 -6256
rect 7148 -6880 7228 -6872
rect 7148 -6934 7158 -6880
rect 7216 -6934 7228 -6880
rect 7148 -6946 7228 -6934
<< via2 >>
rect 6447 -3106 6507 -3102
rect 6447 -3158 6451 -3106
rect 6451 -3158 6503 -3106
rect 6503 -3158 6507 -3106
rect 6447 -3162 6507 -3158
rect 6292 -3514 6358 -3454
rect 7475 -4339 7618 -4188
rect 6580 -4375 6640 -4371
rect 6580 -4427 6584 -4375
rect 6584 -4427 6636 -4375
rect 6636 -4427 6640 -4375
rect 6580 -4431 6640 -4427
<< metal3 >>
rect 6430 -3097 6536 -3084
rect 6430 -3167 6442 -3097
rect 6512 -3167 6536 -3097
rect 6430 -3180 6536 -3167
rect 6286 -3454 6376 -3442
rect 6286 -3514 6292 -3454
rect 6358 -3456 6376 -3454
rect 6358 -3514 6624 -3456
rect 6286 -3516 6624 -3514
rect 6286 -3526 6376 -3516
rect 7433 -4188 7654 -4156
rect 7433 -4339 7475 -4188
rect 7618 -4339 7654 -4188
rect 6549 -4366 6676 -4348
rect 6549 -4436 6575 -4366
rect 6645 -4436 6676 -4366
rect 7433 -4378 7654 -4339
rect 6549 -4459 6676 -4436
<< via3 >>
rect 6442 -3102 6512 -3097
rect 6442 -3162 6447 -3102
rect 6447 -3162 6507 -3102
rect 6507 -3162 6512 -3102
rect 6442 -3167 6512 -3162
rect 7475 -4339 7618 -4188
rect 6575 -4371 6645 -4366
rect 6575 -4431 6580 -4371
rect 6580 -4431 6640 -4371
rect 6640 -4431 6645 -4371
rect 6575 -4436 6645 -4431
<< metal4 >>
rect 8149 -2221 8832 -2093
rect 6441 -3097 6513 -3096
rect 6441 -3167 6442 -3097
rect 6512 -3167 6513 -3097
rect 6441 -3168 6513 -3167
rect 6447 -3228 6510 -3168
rect 6434 -3332 6777 -3228
rect 6436 -3333 6777 -3332
rect 6436 -4371 6496 -3333
rect 7433 -4188 7654 -4156
rect 7433 -4339 7475 -4188
rect 7618 -4196 7654 -4188
rect 8149 -4196 8277 -2221
rect 7618 -4324 8277 -4196
rect 7618 -4339 7654 -4324
rect 6574 -4366 6646 -4365
rect 6574 -4371 6575 -4366
rect 6436 -4431 6575 -4371
rect 6574 -4436 6575 -4431
rect 6645 -4436 6646 -4366
rect 7433 -4378 7654 -4339
rect 6574 -4437 6646 -4436
use bodynmos  bodynmos_1
timestamp 1717180972
transform 1 0 4760 0 1 -5863
box -24 -24 62 52
use bodypmos  bodypmos_0
timestamp 1717180972
transform 1 0 6022 0 1 -2712
box -76 -78 118 110
use sky130_fd_pr__cap_mim_m3_1_FJK8MD  sky130_fd_pr__cap_mim_m3_1_FJK8MD_0
timestamp 1717180972
transform 0 1 6856 -1 0 -3592
box -386 -240 386 240
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_0
timestamp 1717180972
transform 1 0 8010 0 1 -6069
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_1
timestamp 1717180972
transform -1 0 7605 0 1 -6068
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_2
timestamp 1717180972
transform 1 0 7201 0 1 -6068
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_3
timestamp 1717180972
transform -1 0 6795 0 1 -6070
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_4
timestamp 1717180972
transform 1 0 6389 0 1 -6070
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_24PS5X  sky130_fd_pr__nfet_01v8_24PS5X_5
timestamp 1717180972
transform -1 0 5983 0 1 -6070
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_5U3WHE  sky130_fd_pr__pfet_01v8_5U3WHE_0
timestamp 1717180972
transform 1 0 6307 0 1 -2694
box -109 -162 109 162
use sky130_fd_pr__res_xhigh_po_0p35_6R3NZW  sky130_fd_pr__res_xhigh_po_0p35_6R3NZW_0
timestamp 1717180972
transform 1 0 4915 0 1 -6573
box -35 -482 35 482
use sky130_fd_pr__cap_mim_m3_1_F2GAMD  XC8
timestamp 1717180972
transform 1 0 9115 0 1 -5014
box -386 -3240 386 3240
use sky130_fd_pr__pfet_01v8_5U3WHE  XM29
timestamp 1717180972
transform 1 0 6609 0 1 -2694
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_5U3WHE  XM39
timestamp 1717180972
transform -1 0 6219 0 1 -2694
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_5U3WHE  XM42
timestamp 1717180972
transform -1 0 6521 0 1 -2694
box -109 -162 109 162
use sky130_fd_pr__nfet_01v8_WYB6A9  XM43
timestamp 1717180972
transform 1 0 4958 0 1 -5823
box -73 -126 73 126
<< labels >>
rlabel locali 6033 -2552 6059 -2525 1 vdd
port 4 n
rlabel space 4992 -5686 5020 -5659 1 vdd
port 5 n
rlabel metal1 6480 -6928 6506 -6906 1 vref
port 2 n
rlabel metal1 5894 -6751 5921 -6733 1 in1
port 1 n
rlabel locali 5282 -5520 5322 -5494 1 v1
rlabel metal1 5814 -5384 5838 -5354 1 vss
<< end >>
