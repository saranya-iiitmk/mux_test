magic
tech sky130A
magscale 1 2
timestamp 1718685184
<< viali >>
rect 3893 14025 3927 14059
rect 11069 14025 11103 14059
rect 12909 13957 12943 13991
rect 4169 13889 4203 13923
rect 10977 13889 11011 13923
rect 12725 13753 12759 13787
rect 8953 13345 8987 13379
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 8125 13277 8159 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 9689 13277 9723 13311
rect 10241 13277 10275 13311
rect 10517 13209 10551 13243
rect 7481 13141 7515 13175
rect 7941 13141 7975 13175
rect 9873 13141 9907 13175
rect 11989 13141 12023 13175
rect 11621 12937 11655 12971
rect 6545 12869 6579 12903
rect 6745 12869 6779 12903
rect 7021 12869 7055 12903
rect 7757 12869 7791 12903
rect 5641 12801 5675 12835
rect 6101 12801 6135 12835
rect 7205 12801 7239 12835
rect 7481 12801 7515 12835
rect 9781 12801 9815 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 5733 12665 5767 12699
rect 6377 12665 6411 12699
rect 9597 12665 9631 12699
rect 10609 12665 10643 12699
rect 5917 12597 5951 12631
rect 6561 12597 6595 12631
rect 7389 12597 7423 12631
rect 9965 12597 9999 12631
rect 7389 12393 7423 12427
rect 7573 12393 7607 12427
rect 8585 12393 8619 12427
rect 9689 12393 9723 12427
rect 11897 12393 11931 12427
rect 8401 12325 8435 12359
rect 5089 12257 5123 12291
rect 7941 12257 7975 12291
rect 9781 12257 9815 12291
rect 8033 12189 8067 12223
rect 8493 12189 8527 12223
rect 9137 12189 9171 12223
rect 9505 12189 9539 12223
rect 9965 12189 9999 12223
rect 10057 12189 10091 12223
rect 10241 12189 10275 12223
rect 10333 12189 10367 12223
rect 11989 12189 12023 12223
rect 5365 12121 5399 12155
rect 7205 12121 7239 12155
rect 7405 12121 7439 12155
rect 9321 12121 9355 12155
rect 9413 12121 9447 12155
rect 6837 12053 6871 12087
rect 11529 12053 11563 12087
rect 7205 11849 7239 11883
rect 9873 11849 9907 11883
rect 6653 11781 6687 11815
rect 6853 11781 6887 11815
rect 9505 11781 9539 11815
rect 4813 11713 4847 11747
rect 7297 11713 7331 11747
rect 9413 11713 9447 11747
rect 9597 11713 9631 11747
rect 10057 11713 10091 11747
rect 10150 11713 10184 11747
rect 10425 11713 10459 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 12173 11713 12207 11747
rect 11161 11645 11195 11679
rect 11345 11645 11379 11679
rect 11621 11645 11655 11679
rect 7021 11577 7055 11611
rect 9781 11577 9815 11611
rect 4629 11509 4663 11543
rect 6837 11509 6871 11543
rect 9229 11509 9263 11543
rect 10333 11509 10367 11543
rect 11253 11509 11287 11543
rect 11989 11509 12023 11543
rect 12265 11509 12299 11543
rect 4064 11305 4098 11339
rect 6837 11305 6871 11339
rect 8125 11305 8159 11339
rect 9045 11305 9079 11339
rect 11161 11305 11195 11339
rect 3801 11169 3835 11203
rect 6193 11169 6227 11203
rect 7113 11169 7147 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 11713 11169 11747 11203
rect 5825 11101 5859 11135
rect 6101 11101 6135 11135
rect 7021 11101 7055 11135
rect 9229 11101 9263 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 11989 11101 12023 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 8309 11033 8343 11067
rect 8493 11033 8527 11067
rect 6469 10965 6503 10999
rect 11529 10965 11563 10999
rect 4721 10761 4755 10795
rect 6377 10761 6411 10795
rect 10333 10761 10367 10795
rect 10701 10761 10735 10795
rect 11897 10761 11931 10795
rect 6101 10693 6135 10727
rect 6837 10693 6871 10727
rect 8217 10693 8251 10727
rect 8401 10693 8435 10727
rect 9597 10693 9631 10727
rect 4629 10625 4663 10659
rect 5917 10625 5951 10659
rect 6193 10625 6227 10659
rect 7849 10625 7883 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 8493 10625 8527 10659
rect 9781 10625 9815 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 10425 10625 10459 10659
rect 10793 10625 10827 10659
rect 12725 10625 12759 10659
rect 7205 10557 7239 10591
rect 10885 10557 10919 10591
rect 13001 10557 13035 10591
rect 6561 10489 6595 10523
rect 8125 10489 8159 10523
rect 9873 10489 9907 10523
rect 11253 10489 11287 10523
rect 11345 10489 11379 10523
rect 11529 10489 11563 10523
rect 12081 10489 12115 10523
rect 5917 10421 5951 10455
rect 8217 10421 8251 10455
rect 11897 10421 11931 10455
rect 7021 10217 7055 10251
rect 9781 10217 9815 10251
rect 9965 10217 9999 10251
rect 10517 10217 10551 10251
rect 10885 10217 10919 10251
rect 12081 10217 12115 10251
rect 12541 10217 12575 10251
rect 9597 10149 9631 10183
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 6837 10081 6871 10115
rect 7389 10081 7423 10115
rect 12173 10081 12207 10115
rect 3341 10013 3375 10047
rect 7205 10013 7239 10047
rect 9873 10013 9907 10047
rect 10425 10013 10459 10047
rect 11437 10013 11471 10047
rect 11530 10013 11564 10047
rect 11902 10013 11936 10047
rect 12633 10013 12667 10047
rect 9321 9945 9355 9979
rect 11713 9945 11747 9979
rect 11805 9945 11839 9979
rect 3157 9877 3191 9911
rect 10333 9877 10367 9911
rect 6009 9673 6043 9707
rect 9965 9673 9999 9707
rect 11621 9673 11655 9707
rect 2881 9605 2915 9639
rect 4629 9605 4663 9639
rect 8033 9605 8067 9639
rect 12081 9605 12115 9639
rect 4721 9537 4755 9571
rect 5917 9537 5951 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 9689 9537 9723 9571
rect 9781 9537 9815 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11253 9537 11287 9571
rect 11805 9537 11839 9571
rect 2605 9469 2639 9503
rect 9965 9469 9999 9503
rect 11897 9469 11931 9503
rect 9505 9401 9539 9435
rect 10977 9401 11011 9435
rect 4353 9333 4387 9367
rect 7389 9333 7423 9367
rect 10517 9333 10551 9367
rect 11069 9333 11103 9367
rect 12081 9333 12115 9367
rect 7205 9129 7239 9163
rect 8309 9129 8343 9163
rect 12265 9129 12299 9163
rect 4997 9061 5031 9095
rect 3249 8993 3283 9027
rect 5273 8993 5307 9027
rect 7297 8993 7331 9027
rect 7849 8993 7883 9027
rect 3525 8925 3559 8959
rect 4236 8925 4270 8959
rect 4721 8925 4755 8959
rect 5457 8925 5491 8959
rect 8217 8925 8251 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 12357 8925 12391 8959
rect 2973 8857 3007 8891
rect 4445 8857 4479 8891
rect 5733 8857 5767 8891
rect 1501 8789 1535 8823
rect 3433 8789 3467 8823
rect 4077 8789 4111 8823
rect 4353 8789 4387 8823
rect 4813 8789 4847 8823
rect 11437 8789 11471 8823
rect 3249 8585 3283 8619
rect 3341 8585 3375 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 12357 8585 12391 8619
rect 2421 8517 2455 8551
rect 3525 8517 3559 8551
rect 3985 8517 4019 8551
rect 6377 8517 6411 8551
rect 2329 8449 2363 8483
rect 2513 8449 2547 8483
rect 2605 8449 2639 8483
rect 2789 8449 2823 8483
rect 2881 8449 2915 8483
rect 2973 8449 3007 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 5917 8449 5951 8483
rect 6193 8449 6227 8483
rect 12081 8449 12115 8483
rect 12909 8381 12943 8415
rect 3893 8313 3927 8347
rect 3525 8245 3559 8279
rect 7665 8245 7699 8279
rect 12173 8245 12207 8279
rect 2605 8041 2639 8075
rect 3065 8041 3099 8075
rect 5549 8041 5583 8075
rect 12909 8041 12943 8075
rect 2237 7905 2271 7939
rect 11437 7905 11471 7939
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 2789 7837 2823 7871
rect 2973 7837 3007 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 7021 7837 7055 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 9689 7837 9723 7871
rect 11161 7837 11195 7871
rect 8953 7769 8987 7803
rect 9137 7769 9171 7803
rect 2237 7701 2271 7735
rect 8033 7701 8067 7735
rect 8401 7701 8435 7735
rect 9321 7701 9355 7735
rect 9505 7701 9539 7735
rect 2697 7497 2731 7531
rect 5733 7429 5767 7463
rect 8769 7429 8803 7463
rect 9505 7429 9539 7463
rect 11161 7429 11195 7463
rect 2605 7361 2639 7395
rect 2789 7361 2823 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 9056 7361 9090 7395
rect 9229 7361 9263 7395
rect 11253 7361 11287 7395
rect 12173 7361 12207 7395
rect 5365 7225 5399 7259
rect 5917 7225 5951 7259
rect 5733 7157 5767 7191
rect 6009 7157 6043 7191
rect 6653 7157 6687 7191
rect 7297 7157 7331 7191
rect 10977 7157 11011 7191
rect 12265 7157 12299 7191
rect 1672 6953 1706 6987
rect 8401 6953 8435 6987
rect 8585 6953 8619 6987
rect 9137 6953 9171 6987
rect 9321 6953 9355 6987
rect 9965 6953 9999 6987
rect 10609 6953 10643 6987
rect 1409 6817 1443 6851
rect 5549 6817 5583 6851
rect 5825 6817 5859 6851
rect 11161 6817 11195 6851
rect 3433 6749 3467 6783
rect 4905 6749 4939 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 10885 6749 10919 6783
rect 3341 6681 3375 6715
rect 4169 6681 4203 6715
rect 4353 6681 4387 6715
rect 5089 6681 5123 6715
rect 5273 6681 5307 6715
rect 5457 6681 5491 6715
rect 9321 6681 9355 6715
rect 10149 6681 10183 6715
rect 11437 6681 11471 6715
rect 3157 6613 3191 6647
rect 4537 6613 4571 6647
rect 4721 6613 4755 6647
rect 7297 6613 7331 6647
rect 8401 6613 8435 6647
rect 9781 6613 9815 6647
rect 9939 6613 9973 6647
rect 10609 6613 10643 6647
rect 10793 6613 10827 6647
rect 11069 6613 11103 6647
rect 12909 6613 12943 6647
rect 3893 6409 3927 6443
rect 8585 6409 8619 6443
rect 9505 6409 9539 6443
rect 9873 6409 9907 6443
rect 10333 6409 10367 6443
rect 4045 6341 4079 6375
rect 4261 6341 4295 6375
rect 4629 6341 4663 6375
rect 8217 6341 8251 6375
rect 9689 6341 9723 6375
rect 9965 6341 9999 6375
rect 10149 6341 10183 6375
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3525 6273 3559 6307
rect 8401 6273 8435 6307
rect 9597 6273 9631 6307
rect 12725 6273 12759 6307
rect 3341 6205 3375 6239
rect 4360 6205 4394 6239
rect 6101 6205 6135 6239
rect 9321 6205 9355 6239
rect 13001 6205 13035 6239
rect 2421 6069 2455 6103
rect 2789 6069 2823 6103
rect 3709 6069 3743 6103
rect 4077 6069 4111 6103
rect 4353 5865 4387 5899
rect 4537 5865 4571 5899
rect 6469 5865 6503 5899
rect 7959 5865 7993 5899
rect 1501 5729 1535 5763
rect 1777 5729 1811 5763
rect 3985 5729 4019 5763
rect 4629 5729 4663 5763
rect 8217 5729 8251 5763
rect 6377 5661 6411 5695
rect 8309 5661 8343 5695
rect 4353 5593 4387 5627
rect 8401 5593 8435 5627
rect 3249 5525 3283 5559
rect 2789 5321 2823 5355
rect 4997 5321 5031 5355
rect 5365 5321 5399 5355
rect 5733 5321 5767 5355
rect 8769 5321 8803 5355
rect 11177 5321 11211 5355
rect 11345 5321 11379 5355
rect 2973 5253 3007 5287
rect 3801 5253 3835 5287
rect 4169 5253 4203 5287
rect 5181 5253 5215 5287
rect 5549 5253 5583 5287
rect 8283 5253 8317 5287
rect 8401 5253 8435 5287
rect 10517 5253 10551 5287
rect 10977 5253 11011 5287
rect 2145 5185 2179 5219
rect 3341 5185 3375 5219
rect 3985 5185 4019 5219
rect 5273 5185 5307 5219
rect 5825 5185 5859 5219
rect 7481 5185 7515 5219
rect 8493 5185 8527 5219
rect 8585 5185 8619 5219
rect 9321 5185 9355 5219
rect 9781 5185 9815 5219
rect 10241 5185 10275 5219
rect 10425 5185 10459 5219
rect 10701 5185 10735 5219
rect 11713 5185 11747 5219
rect 12173 5185 12207 5219
rect 2421 5117 2455 5151
rect 8033 5117 8067 5151
rect 8125 5117 8159 5151
rect 10333 5117 10367 5151
rect 2973 4981 3007 5015
rect 9229 4981 9263 5015
rect 9689 4981 9723 5015
rect 10885 4981 10919 5015
rect 11161 4981 11195 5015
rect 11529 4981 11563 5015
rect 12265 4981 12299 5015
rect 10701 4777 10735 4811
rect 2973 4641 3007 4675
rect 11437 4641 11471 4675
rect 1409 4573 1443 4607
rect 2697 4573 2731 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 1593 4437 1627 4471
rect 12909 4437 12943 4471
rect 8585 4233 8619 4267
rect 10241 4233 10275 4267
rect 10977 4233 11011 4267
rect 5641 4165 5675 4199
rect 11161 4165 11195 4199
rect 2237 4097 2271 4131
rect 2881 4097 2915 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 7665 4097 7699 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 8861 4097 8895 4131
rect 9413 4097 9447 4131
rect 10391 4097 10425 4131
rect 10885 4097 10919 4131
rect 11713 4097 11747 4131
rect 12357 4097 12391 4131
rect 12909 4097 12943 4131
rect 3709 4029 3743 4063
rect 5825 4029 5859 4063
rect 6009 4029 6043 4063
rect 6745 4029 6779 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 11621 4029 11655 4063
rect 2605 3961 2639 3995
rect 4077 3961 4111 3995
rect 5273 3961 5307 3995
rect 7021 3961 7055 3995
rect 7113 3961 7147 3995
rect 7941 3961 7975 3995
rect 11161 3961 11195 3995
rect 2697 3893 2731 3927
rect 2973 3893 3007 3927
rect 3341 3893 3375 3927
rect 4169 3893 4203 3927
rect 4629 3893 4663 3927
rect 5181 3893 5215 3927
rect 5917 3893 5951 3927
rect 8861 3893 8895 3927
rect 9137 3893 9171 3927
rect 9321 3893 9355 3927
rect 12081 3893 12115 3927
rect 1685 3689 1719 3723
rect 2329 3689 2363 3723
rect 2697 3689 2731 3723
rect 4537 3689 4571 3723
rect 5549 3689 5583 3723
rect 7021 3689 7055 3723
rect 7389 3689 7423 3723
rect 8953 3689 8987 3723
rect 9413 3689 9447 3723
rect 10241 3689 10275 3723
rect 10977 3689 11011 3723
rect 12909 3689 12943 3723
rect 1961 3621 1995 3655
rect 2513 3621 2547 3655
rect 3525 3621 3559 3655
rect 5733 3621 5767 3655
rect 6377 3621 6411 3655
rect 4077 3553 4111 3587
rect 4169 3553 4203 3587
rect 5917 3553 5951 3587
rect 7113 3553 7147 3587
rect 8033 3553 8067 3587
rect 8125 3553 8159 3587
rect 10517 3553 10551 3587
rect 11161 3553 11195 3587
rect 1409 3485 1443 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4353 3485 4387 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 5825 3485 5859 3519
rect 6101 3485 6135 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 7205 3485 7239 3519
rect 7606 3485 7640 3519
rect 8401 3485 8435 3519
rect 8769 3485 8803 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 9505 3485 9539 3519
rect 9597 3485 9631 3519
rect 9690 3485 9724 3519
rect 9965 3485 9999 3519
rect 10062 3485 10096 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 10885 3485 10919 3519
rect 2973 3417 3007 3451
rect 6929 3417 6963 3451
rect 8493 3417 8527 3451
rect 8585 3417 8619 3451
rect 9873 3417 9907 3451
rect 11437 3417 11471 3451
rect 1869 3349 1903 3383
rect 2329 3349 2363 3383
rect 2881 3349 2915 3383
rect 3341 3349 3375 3383
rect 7481 3349 7515 3383
rect 7665 3349 7699 3383
rect 8217 3349 8251 3383
rect 2973 3145 3007 3179
rect 3065 3145 3099 3179
rect 4445 3145 4479 3179
rect 5641 3145 5675 3179
rect 6929 3145 6963 3179
rect 7297 3145 7331 3179
rect 7941 3145 7975 3179
rect 8769 3145 8803 3179
rect 9689 3145 9723 3179
rect 12265 3145 12299 3179
rect 12541 3145 12575 3179
rect 4077 3077 4111 3111
rect 5365 3077 5399 3111
rect 5733 3077 5767 3111
rect 7573 3077 7607 3111
rect 8493 3077 8527 3111
rect 2513 3009 2547 3043
rect 3525 3009 3559 3043
rect 3893 3009 3927 3043
rect 3985 3009 4019 3043
rect 4261 3009 4295 3043
rect 4353 3009 4387 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5457 3009 5491 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 6469 3009 6503 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 7757 3009 7791 3043
rect 8263 3009 8297 3043
rect 8401 3009 8435 3043
rect 8585 3009 8619 3043
rect 9137 3009 9171 3043
rect 9413 3009 9447 3043
rect 9505 3009 9539 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 12449 3009 12483 3043
rect 13001 3009 13035 3043
rect 4905 2941 4939 2975
rect 6653 2941 6687 2975
rect 9229 2941 9263 2975
rect 4537 2873 4571 2907
rect 12817 2873 12851 2907
rect 2789 2805 2823 2839
rect 3433 2805 3467 2839
rect 3709 2805 3743 2839
rect 6469 2805 6503 2839
rect 1593 2601 1627 2635
rect 2789 2601 2823 2635
rect 4353 2601 4387 2635
rect 5917 2601 5951 2635
rect 8953 2601 8987 2635
rect 10425 2601 10459 2635
rect 12817 2601 12851 2635
rect 7297 2533 7331 2567
rect 11805 2465 11839 2499
rect 1409 2397 1443 2431
rect 2605 2397 2639 2431
rect 4169 2397 4203 2431
rect 5733 2397 5767 2431
rect 6745 2397 6779 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 11529 2397 11563 2431
rect 12909 2329 12943 2363
<< metal1 >>
rect 1104 14170 13499 14192
rect 1104 14118 4008 14170
rect 4060 14118 4072 14170
rect 4124 14118 4136 14170
rect 4188 14118 4200 14170
rect 4252 14118 4264 14170
rect 4316 14118 7067 14170
rect 7119 14118 7131 14170
rect 7183 14118 7195 14170
rect 7247 14118 7259 14170
rect 7311 14118 7323 14170
rect 7375 14118 10126 14170
rect 10178 14118 10190 14170
rect 10242 14118 10254 14170
rect 10306 14118 10318 14170
rect 10370 14118 10382 14170
rect 10434 14118 13185 14170
rect 13237 14118 13249 14170
rect 13301 14118 13313 14170
rect 13365 14118 13377 14170
rect 13429 14118 13441 14170
rect 13493 14118 13499 14170
rect 1104 14096 13499 14118
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 3660 14028 3893 14056
rect 3660 14016 3666 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10836 14028 11069 14056
rect 10836 14016 10842 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 12897 13991 12955 13997
rect 12897 13957 12909 13991
rect 12943 13988 12955 13991
rect 13262 13988 13268 14000
rect 12943 13960 13268 13988
rect 12943 13957 12955 13960
rect 12897 13951 12955 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 6270 13920 6276 13932
rect 4203 13892 6276 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 12710 13744 12716 13796
rect 12768 13744 12774 13796
rect 1104 13626 13340 13648
rect 1104 13574 2479 13626
rect 2531 13574 2543 13626
rect 2595 13574 2607 13626
rect 2659 13574 2671 13626
rect 2723 13574 2735 13626
rect 2787 13574 5538 13626
rect 5590 13574 5602 13626
rect 5654 13574 5666 13626
rect 5718 13574 5730 13626
rect 5782 13574 5794 13626
rect 5846 13574 8597 13626
rect 8649 13574 8661 13626
rect 8713 13574 8725 13626
rect 8777 13574 8789 13626
rect 8841 13574 8853 13626
rect 8905 13574 11656 13626
rect 11708 13574 11720 13626
rect 11772 13574 11784 13626
rect 11836 13574 11848 13626
rect 11900 13574 11912 13626
rect 11964 13574 13340 13626
rect 1104 13552 13340 13574
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 6788 13348 8953 13376
rect 6788 13336 6794 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 6972 13280 7297 13308
rect 6972 13268 6978 13280
rect 7285 13277 7297 13280
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 7515 13280 7788 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 7760 13184 7788 13280
rect 8110 13268 8116 13320
rect 8168 13268 8174 13320
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9355 13280 9689 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9824 13280 10241 13308
rect 9824 13268 9830 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 10505 13243 10563 13249
rect 10505 13240 10517 13243
rect 9876 13212 10517 13240
rect 7466 13132 7472 13184
rect 7524 13132 7530 13184
rect 7742 13132 7748 13184
rect 7800 13132 7806 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 9876 13181 9904 13212
rect 10505 13209 10517 13212
rect 10551 13209 10563 13243
rect 10505 13203 10563 13209
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7892 13144 7941 13172
rect 7892 13132 7898 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 9861 13175 9919 13181
rect 9861 13141 9873 13175
rect 9907 13141 9919 13175
rect 9861 13135 9919 13141
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 1104 13082 13499 13104
rect 1104 13030 4008 13082
rect 4060 13030 4072 13082
rect 4124 13030 4136 13082
rect 4188 13030 4200 13082
rect 4252 13030 4264 13082
rect 4316 13030 7067 13082
rect 7119 13030 7131 13082
rect 7183 13030 7195 13082
rect 7247 13030 7259 13082
rect 7311 13030 7323 13082
rect 7375 13030 10126 13082
rect 10178 13030 10190 13082
rect 10242 13030 10254 13082
rect 10306 13030 10318 13082
rect 10370 13030 10382 13082
rect 10434 13030 13185 13082
rect 13237 13030 13249 13082
rect 13301 13030 13313 13082
rect 13365 13030 13377 13082
rect 13429 13030 13441 13082
rect 13493 13030 13499 13082
rect 1104 13008 13499 13030
rect 9766 12968 9772 12980
rect 7484 12940 9772 12968
rect 6533 12903 6591 12909
rect 6533 12869 6545 12903
rect 6579 12900 6591 12903
rect 6638 12900 6644 12912
rect 6579 12872 6644 12900
rect 6579 12869 6591 12872
rect 6533 12863 6591 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6730 12860 6736 12912
rect 6788 12860 6794 12912
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7009 12903 7067 12909
rect 7009 12900 7021 12903
rect 6972 12872 7021 12900
rect 6972 12860 6978 12872
rect 7009 12869 7021 12872
rect 7055 12869 7067 12903
rect 7009 12863 7067 12869
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 6089 12835 6147 12841
rect 5675 12804 5709 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 7193 12835 7251 12841
rect 6135 12804 6408 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5644 12764 5672 12795
rect 5500 12736 6132 12764
rect 5500 12724 5506 12736
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 5767 12668 6040 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 6012 12640 6040 12668
rect 5902 12588 5908 12640
rect 5960 12588 5966 12640
rect 5994 12588 6000 12640
rect 6052 12588 6058 12640
rect 6104 12628 6132 12736
rect 6380 12705 6408 12804
rect 7193 12801 7205 12835
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7208 12764 7236 12795
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7484 12841 7512 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11606 12928 11612 12980
rect 11664 12928 11670 12980
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 7834 12900 7840 12912
rect 7791 12872 7840 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 7834 12860 7840 12872
rect 7892 12860 7898 12912
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 12710 12900 12716 12912
rect 10704 12872 12716 12900
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7340 12804 7481 12832
rect 7340 12792 7346 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 10704 12841 10732 12872
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 10836 12804 11713 12832
rect 10836 12792 10842 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 7742 12764 7748 12776
rect 7208 12736 7748 12764
rect 7742 12724 7748 12736
rect 7800 12764 7806 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 7800 12736 9229 12764
rect 7800 12724 7806 12736
rect 9217 12733 9229 12736
rect 9263 12764 9275 12767
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9263 12736 9505 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9493 12733 9505 12736
rect 9539 12764 9551 12767
rect 9858 12764 9864 12776
rect 9539 12736 9864 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12665 6423 12699
rect 9585 12699 9643 12705
rect 6365 12659 6423 12665
rect 6472 12668 7512 12696
rect 6472 12628 6500 12668
rect 6104 12600 6500 12628
rect 6546 12588 6552 12640
rect 6604 12588 6610 12640
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 7484 12628 7512 12668
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10042 12696 10048 12708
rect 9631 12668 10048 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10042 12656 10048 12668
rect 10100 12696 10106 12708
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10100 12668 10609 12696
rect 10100 12656 10106 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 8202 12628 8208 12640
rect 7484 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9953 12631 10011 12637
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10134 12628 10140 12640
rect 9999 12600 10140 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 1104 12538 13340 12560
rect 1104 12486 2479 12538
rect 2531 12486 2543 12538
rect 2595 12486 2607 12538
rect 2659 12486 2671 12538
rect 2723 12486 2735 12538
rect 2787 12486 5538 12538
rect 5590 12486 5602 12538
rect 5654 12486 5666 12538
rect 5718 12486 5730 12538
rect 5782 12486 5794 12538
rect 5846 12486 8597 12538
rect 8649 12486 8661 12538
rect 8713 12486 8725 12538
rect 8777 12486 8789 12538
rect 8841 12486 8853 12538
rect 8905 12486 11656 12538
rect 11708 12486 11720 12538
rect 11772 12486 11784 12538
rect 11836 12486 11848 12538
rect 11900 12486 11912 12538
rect 11964 12486 13340 12538
rect 1104 12464 13340 12486
rect 7282 12424 7288 12436
rect 5184 12396 7288 12424
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 5184 12288 5212 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 7466 12424 7472 12436
rect 7423 12396 7472 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 7561 12427 7619 12433
rect 7561 12393 7573 12427
rect 7607 12424 7619 12427
rect 8110 12424 8116 12436
rect 7607 12396 8116 12424
rect 7607 12393 7619 12396
rect 7561 12387 7619 12393
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8536 12396 8585 12424
rect 8536 12384 8542 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9122 12384 9128 12436
rect 9180 12384 9186 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9766 12424 9772 12436
rect 9723 12396 9772 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10778 12424 10784 12436
rect 9876 12396 10784 12424
rect 7374 12288 7380 12300
rect 5132 12260 5212 12288
rect 7300 12260 7380 12288
rect 5132 12248 5138 12260
rect 5353 12155 5411 12161
rect 5353 12121 5365 12155
rect 5399 12152 5411 12155
rect 5626 12152 5632 12164
rect 5399 12124 5632 12152
rect 5399 12121 5411 12124
rect 5353 12115 5411 12121
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 5994 12112 6000 12164
rect 6052 12112 6058 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6788 12124 7205 12152
rect 6788 12112 6794 12124
rect 7193 12121 7205 12124
rect 7239 12121 7251 12155
rect 7300 12152 7328 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7484 12288 7512 12384
rect 8389 12359 8447 12365
rect 8389 12325 8401 12359
rect 8435 12356 8447 12359
rect 9140 12356 9168 12384
rect 9876 12356 9904 12396
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11026 12396 11897 12424
rect 10042 12356 10048 12368
rect 8435 12328 9168 12356
rect 9232 12328 9904 12356
rect 9968 12328 10048 12356
rect 8435 12325 8447 12328
rect 8389 12319 8447 12325
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7484 12260 7941 12288
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 9232 12288 9260 12328
rect 8260 12260 9260 12288
rect 8260 12248 8266 12260
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8496 12229 8524 12260
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 9732 12260 9781 12288
rect 9732 12248 9738 12260
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 9968 12229 9996 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10134 12316 10140 12368
rect 10192 12316 10198 12368
rect 10226 12316 10232 12368
rect 10284 12356 10290 12368
rect 10284 12328 10364 12356
rect 10284 12316 10290 12328
rect 10152 12288 10180 12316
rect 10336 12288 10364 12328
rect 11026 12288 11054 12396
rect 11885 12393 11897 12396
rect 11931 12424 11943 12427
rect 11974 12424 11980 12436
rect 11931 12396 11980 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12710 12288 12716 12300
rect 10152 12260 10272 12288
rect 10244 12229 10272 12260
rect 10336 12260 11054 12288
rect 11992 12260 12716 12288
rect 10336 12229 10364 12260
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 7393 12155 7451 12161
rect 7393 12152 7405 12155
rect 7300 12124 7405 12152
rect 7193 12115 7251 12121
rect 7393 12121 7405 12124
rect 7439 12121 7451 12155
rect 7393 12115 7451 12121
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 6362 12084 6368 12096
rect 4120 12056 6368 12084
rect 4120 12044 4126 12056
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 6822 12044 6828 12096
rect 6880 12044 6886 12096
rect 7208 12084 7236 12115
rect 9306 12112 9312 12164
rect 9364 12112 9370 12164
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 7558 12084 7564 12096
rect 7208 12056 7564 12084
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 9416 12084 9444 12115
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10060 12152 10088 12183
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11992 12229 12020 12260
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11480 12192 11989 12220
rect 11480 12180 11486 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 9916 12124 10088 12152
rect 9916 12112 9922 12124
rect 9950 12084 9956 12096
rect 9416 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10060 12084 10088 12124
rect 10502 12084 10508 12096
rect 10060 12056 10508 12084
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11514 12044 11520 12096
rect 11572 12044 11578 12096
rect 1104 11994 13499 12016
rect 1104 11942 4008 11994
rect 4060 11942 4072 11994
rect 4124 11942 4136 11994
rect 4188 11942 4200 11994
rect 4252 11942 4264 11994
rect 4316 11942 7067 11994
rect 7119 11942 7131 11994
rect 7183 11942 7195 11994
rect 7247 11942 7259 11994
rect 7311 11942 7323 11994
rect 7375 11942 10126 11994
rect 10178 11942 10190 11994
rect 10242 11942 10254 11994
rect 10306 11942 10318 11994
rect 10370 11942 10382 11994
rect 10434 11942 13185 11994
rect 13237 11942 13249 11994
rect 13301 11942 13313 11994
rect 13365 11942 13377 11994
rect 13429 11942 13441 11994
rect 13493 11942 13499 11994
rect 1104 11920 13499 11942
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6604 11852 7205 11880
rect 6604 11840 6610 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9180 11852 9873 11880
rect 9180 11840 9186 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10042 11840 10048 11892
rect 10100 11840 10106 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11781 6699 11815
rect 6641 11775 6699 11781
rect 6841 11815 6899 11821
rect 6841 11781 6853 11815
rect 6887 11812 6899 11815
rect 9493 11815 9551 11821
rect 6887 11784 7052 11812
rect 6887 11781 6899 11784
rect 6841 11775 6899 11781
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5902 11744 5908 11756
rect 4847 11716 5908 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 6656 11676 6684 11775
rect 7024 11756 7052 11784
rect 9493 11781 9505 11815
rect 9539 11812 9551 11815
rect 10060 11812 10088 11840
rect 9539 11784 10088 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 7006 11704 7012 11756
rect 7064 11704 7070 11756
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 6822 11676 6828 11688
rect 6656 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7300 11676 7328 11707
rect 6972 11648 7328 11676
rect 9416 11676 9444 11707
rect 9582 11704 9588 11756
rect 9640 11704 9646 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 9490 11676 9496 11688
rect 9416 11648 9496 11676
rect 6972 11636 6978 11648
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 10060 11676 10088 11707
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10192 11716 10237 11744
rect 10192 11704 10198 11716
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10376 11716 10425 11744
rect 10376 11704 10382 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10560 11716 11069 11744
rect 10560 11704 10566 11716
rect 11057 11713 11069 11716
rect 11103 11744 11115 11747
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11103 11716 11713 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11992 11744 12020 11840
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11992 11716 12173 11744
rect 11701 11707 11759 11713
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 11146 11676 11152 11688
rect 9548 11648 11152 11676
rect 9548 11636 9554 11648
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 11514 11676 11520 11688
rect 11379 11648 11520 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 6932 11608 6960 11636
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6932 11580 7021 11608
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 7009 11571 7067 11577
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 9824 11580 10364 11608
rect 9824 11568 9830 11580
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7190 11540 7196 11552
rect 6871 11512 7196 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8076 11512 9229 11540
rect 8076 11500 8082 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9217 11503 9275 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10226 11540 10232 11552
rect 9456 11512 10232 11540
rect 9456 11500 9462 11512
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10336 11549 10364 11580
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10686 11540 10692 11552
rect 10367 11512 10692 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11238 11500 11244 11552
rect 11296 11500 11302 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11624 11540 11652 11639
rect 11388 11512 11652 11540
rect 11388 11500 11394 11512
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12250 11500 12256 11552
rect 12308 11500 12314 11552
rect 1104 11450 13340 11472
rect 1104 11398 2479 11450
rect 2531 11398 2543 11450
rect 2595 11398 2607 11450
rect 2659 11398 2671 11450
rect 2723 11398 2735 11450
rect 2787 11398 5538 11450
rect 5590 11398 5602 11450
rect 5654 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 8597 11450
rect 8649 11398 8661 11450
rect 8713 11398 8725 11450
rect 8777 11398 8789 11450
rect 8841 11398 8853 11450
rect 8905 11398 11656 11450
rect 11708 11398 11720 11450
rect 11772 11398 11784 11450
rect 11836 11398 11848 11450
rect 11900 11398 11912 11450
rect 11964 11398 13340 11450
rect 1104 11376 13340 11398
rect 4052 11339 4110 11345
rect 4052 11305 4064 11339
rect 4098 11336 4110 11339
rect 4614 11336 4620 11348
rect 4098 11308 4620 11336
rect 4098 11305 4110 11308
rect 4052 11299 4110 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6696 11308 6837 11336
rect 6696 11296 6702 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 6972 11308 7328 11336
rect 6972 11296 6978 11308
rect 7006 11268 7012 11280
rect 6196 11240 7012 11268
rect 6196 11212 6224 11240
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7300 11268 7328 11308
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7616 11308 8125 11336
rect 7616 11296 7622 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8113 11299 8171 11305
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9306 11336 9312 11348
rect 9079 11308 9312 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9950 11296 9956 11348
rect 10008 11336 10014 11348
rect 11054 11336 11060 11348
rect 10008 11308 11060 11336
rect 10008 11296 10014 11308
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11146 11296 11152 11348
rect 11204 11296 11210 11348
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 9968 11268 9996 11296
rect 11440 11268 11468 11296
rect 7300 11240 9996 11268
rect 11026 11240 11928 11268
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 3835 11172 5120 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 5092 11144 5120 11172
rect 6178 11160 6184 11212
rect 6236 11160 6242 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6932 11172 7113 11200
rect 6932 11144 6960 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7300 11209 7328 11240
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 9766 11200 9772 11212
rect 7285 11163 7343 11169
rect 9232 11172 9772 11200
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 5859 11104 6101 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 6104 11064 6132 11095
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7742 11132 7748 11144
rect 7055 11104 7748 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 9232 11141 9260 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11026 11200 11054 11240
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10928 11172 11054 11200
rect 11164 11172 11713 11200
rect 10928 11160 10934 11172
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9398 11132 9404 11144
rect 9355 11104 9404 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 6104 11036 7236 11064
rect 7208 11008 7236 11036
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 8297 11067 8355 11073
rect 8297 11064 8309 11067
rect 8076 11036 8309 11064
rect 8076 11024 8082 11036
rect 8297 11033 8309 11036
rect 8343 11033 8355 11067
rect 8297 11027 8355 11033
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 8444 11036 8493 11064
rect 8444 11024 8450 11036
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8481 11027 8539 11033
rect 6457 10999 6515 11005
rect 6457 10965 6469 10999
rect 6503 10996 6515 10999
rect 6638 10996 6644 11008
rect 6503 10968 6644 10996
rect 6503 10965 6515 10968
rect 6457 10959 6515 10965
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 9324 10996 9352 11095
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 10502 11132 10508 11144
rect 9631 11104 10508 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 11164 11132 11192 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11026 11104 11192 11132
rect 11241 11135 11299 11141
rect 11026 11064 11054 11104
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 11330 11132 11336 11144
rect 11287 11104 11336 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 10060 11036 11054 11064
rect 10060 11008 10088 11036
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11256 11064 11284 11095
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 11514 11132 11520 11144
rect 11471 11104 11520 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 11204 11036 11284 11064
rect 11900 11064 11928 11240
rect 11992 11172 12296 11200
rect 11992 11141 12020 11172
rect 12268 11144 12296 11172
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12084 11064 12112 11095
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 11900 11036 12112 11064
rect 11204 11024 11210 11036
rect 7248 10968 9352 10996
rect 7248 10956 7254 10968
rect 10042 10956 10048 11008
rect 10100 10956 10106 11008
rect 11514 10956 11520 11008
rect 11572 10956 11578 11008
rect 1104 10906 13499 10928
rect 1104 10854 4008 10906
rect 4060 10854 4072 10906
rect 4124 10854 4136 10906
rect 4188 10854 4200 10906
rect 4252 10854 4264 10906
rect 4316 10854 7067 10906
rect 7119 10854 7131 10906
rect 7183 10854 7195 10906
rect 7247 10854 7259 10906
rect 7311 10854 7323 10906
rect 7375 10854 10126 10906
rect 10178 10854 10190 10906
rect 10242 10854 10254 10906
rect 10306 10854 10318 10906
rect 10370 10854 10382 10906
rect 10434 10854 13185 10906
rect 13237 10854 13249 10906
rect 13301 10854 13313 10906
rect 13365 10854 13377 10906
rect 13429 10854 13441 10906
rect 13493 10854 13499 10906
rect 1104 10832 13499 10854
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 5442 10752 5448 10804
rect 5500 10752 5506 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 5960 10764 6377 10792
rect 5960 10752 5966 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 6472 10764 8340 10792
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 5460 10656 5488 10752
rect 6089 10727 6147 10733
rect 6089 10693 6101 10727
rect 6135 10724 6147 10727
rect 6472 10724 6500 10764
rect 6135 10696 6500 10724
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6696 10696 6837 10724
rect 6696 10684 6702 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 6825 10687 6883 10693
rect 8036 10696 8217 10724
rect 8036 10668 8064 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 4663 10628 5488 10656
rect 5905 10659 5963 10665
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 5920 10588 5948 10619
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 7006 10656 7012 10668
rect 6236 10628 7012 10656
rect 6236 10616 6242 10628
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7883 10628 7941 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 5920 10560 7052 10588
rect 6549 10523 6607 10529
rect 6549 10489 6561 10523
rect 6595 10520 6607 10523
rect 6730 10520 6736 10532
rect 6595 10492 6736 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 7024 10520 7052 10560
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 7156 10560 7205 10588
rect 7156 10548 7162 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7760 10588 7788 10616
rect 8128 10588 8156 10619
rect 7760 10560 8156 10588
rect 8312 10588 8340 10764
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 9548 10764 10333 10792
rect 9548 10752 9554 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 10686 10752 10692 10804
rect 10744 10752 10750 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11885 10795 11943 10801
rect 11204 10764 11744 10792
rect 11204 10752 11210 10764
rect 8386 10684 8392 10736
rect 8444 10724 8450 10736
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 8444 10696 9597 10724
rect 8444 10684 8450 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 9674 10684 9680 10736
rect 9732 10684 9738 10736
rect 9968 10696 11560 10724
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 9692 10656 9720 10684
rect 8527 10628 9720 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 9766 10616 9772 10668
rect 9824 10616 9830 10668
rect 9968 10665 9996 10696
rect 11532 10668 11560 10696
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10060 10588 10088 10616
rect 8312 10560 10088 10588
rect 7193 10551 7251 10557
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10428 10588 10456 10619
rect 10192 10560 10456 10588
rect 10192 10548 10198 10560
rect 8113 10523 8171 10529
rect 8113 10520 8125 10523
rect 7024 10492 8125 10520
rect 8113 10489 8125 10492
rect 8159 10489 8171 10523
rect 8113 10483 8171 10489
rect 9861 10523 9919 10529
rect 9861 10489 9873 10523
rect 9907 10520 9919 10523
rect 10594 10520 10600 10532
rect 9907 10492 10600 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10796 10520 10824 10619
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 11716 10656 11744 10764
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 11716 10628 12725 10656
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 10873 10591 10931 10597
rect 10873 10557 10885 10591
rect 10919 10588 10931 10591
rect 11054 10588 11060 10600
rect 10919 10560 11060 10588
rect 10919 10557 10931 10560
rect 10873 10551 10931 10557
rect 11054 10548 11060 10560
rect 11112 10588 11118 10600
rect 12618 10588 12624 10600
rect 11112 10560 12624 10588
rect 11112 10548 11118 10560
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 12986 10548 12992 10600
rect 13044 10548 13050 10600
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 10796 10492 11253 10520
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 11333 10523 11391 10529
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 11514 10520 11520 10532
rect 11379 10492 11520 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 5902 10412 5908 10464
rect 5960 10412 5966 10464
rect 8202 10412 8208 10464
rect 8260 10412 8266 10464
rect 11256 10452 11284 10483
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 11790 10480 11796 10532
rect 11848 10520 11854 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 11848 10492 12081 10520
rect 11848 10480 11854 10492
rect 12069 10489 12081 10492
rect 12115 10520 12127 10523
rect 12250 10520 12256 10532
rect 12115 10492 12256 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 11422 10452 11428 10464
rect 11256 10424 11428 10452
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 11974 10452 11980 10464
rect 11931 10424 11980 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 13340 10384
rect 1104 10310 2479 10362
rect 2531 10310 2543 10362
rect 2595 10310 2607 10362
rect 2659 10310 2671 10362
rect 2723 10310 2735 10362
rect 2787 10310 5538 10362
rect 5590 10310 5602 10362
rect 5654 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 8597 10362
rect 8649 10310 8661 10362
rect 8713 10310 8725 10362
rect 8777 10310 8789 10362
rect 8841 10310 8853 10362
rect 8905 10310 11656 10362
rect 11708 10310 11720 10362
rect 11772 10310 11784 10362
rect 11836 10310 11848 10362
rect 11900 10310 11912 10362
rect 11964 10310 13340 10362
rect 1104 10288 13340 10310
rect 7006 10208 7012 10260
rect 7064 10208 7070 10260
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 9456 10220 9628 10248
rect 9456 10208 9462 10220
rect 9600 10189 9628 10220
rect 9766 10208 9772 10260
rect 9824 10208 9830 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10217 10011 10251
rect 9953 10211 10011 10217
rect 9585 10183 9643 10189
rect 9585 10149 9597 10183
rect 9631 10180 9643 10183
rect 9968 10180 9996 10211
rect 10502 10208 10508 10260
rect 10560 10208 10566 10260
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10652 10220 10885 10248
rect 10652 10208 10658 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 11514 10208 11520 10260
rect 11572 10208 11578 10260
rect 11974 10208 11980 10260
rect 12032 10208 12038 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12158 10248 12164 10260
rect 12115 10220 12164 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12710 10248 12716 10260
rect 12575 10220 12716 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 9631 10152 9996 10180
rect 9631 10149 9643 10152
rect 9585 10143 9643 10149
rect 5074 10072 5080 10124
rect 5132 10072 5138 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5902 10112 5908 10124
rect 5399 10084 5908 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7098 10112 7104 10124
rect 6871 10084 7104 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7098 10072 7104 10084
rect 7156 10112 7162 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 7156 10084 7389 10112
rect 7156 10072 7162 10084
rect 7377 10081 7389 10084
rect 7423 10112 7435 10115
rect 10520 10112 10548 10208
rect 7423 10084 10548 10112
rect 11532 10112 11560 10208
rect 11992 10112 12020 10208
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 11532 10084 11744 10112
rect 11992 10084 12173 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 9861 10047 9919 10053
rect 7239 10016 7788 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 5994 9936 6000 9988
rect 6052 9936 6058 9988
rect 7760 9920 7788 10016
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9861 10007 9919 10013
rect 10336 10016 10425 10044
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 9876 9976 9904 10007
rect 10042 9976 10048 9988
rect 9355 9948 10048 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 10042 9936 10048 9948
rect 10100 9936 10106 9988
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10336 9917 10364 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11296 10016 11437 10044
rect 11296 10004 11302 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11716 10044 11744 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 11890 10047 11948 10053
rect 11890 10044 11902 10047
rect 11716 10016 11902 10044
rect 11890 10013 11902 10016
rect 11936 10013 11948 10047
rect 11890 10007 11948 10013
rect 12066 10004 12072 10056
rect 12124 10004 12130 10056
rect 12250 10004 12256 10056
rect 12308 10004 12314 10056
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9945 11759 9979
rect 11701 9939 11759 9945
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9976 11851 9979
rect 12084 9976 12112 10004
rect 11839 9948 12112 9976
rect 11839 9945 11851 9948
rect 11793 9939 11851 9945
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10008 9880 10333 9908
rect 10008 9868 10014 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 11716 9908 11744 9939
rect 12268 9908 12296 10004
rect 11716 9880 12296 9908
rect 10321 9871 10379 9877
rect 1104 9818 13499 9840
rect 1104 9766 4008 9818
rect 4060 9766 4072 9818
rect 4124 9766 4136 9818
rect 4188 9766 4200 9818
rect 4252 9766 4264 9818
rect 4316 9766 7067 9818
rect 7119 9766 7131 9818
rect 7183 9766 7195 9818
rect 7247 9766 7259 9818
rect 7311 9766 7323 9818
rect 7375 9766 10126 9818
rect 10178 9766 10190 9818
rect 10242 9766 10254 9818
rect 10306 9766 10318 9818
rect 10370 9766 10382 9818
rect 10434 9766 13185 9818
rect 13237 9766 13249 9818
rect 13301 9766 13313 9818
rect 13365 9766 13377 9818
rect 13429 9766 13441 9818
rect 13493 9766 13499 9818
rect 1104 9744 13499 9766
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 5500 9676 5948 9704
rect 5500 9664 5506 9676
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3142 9636 3148 9648
rect 2915 9608 3148 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4094 9608 4629 9636
rect 4617 9605 4629 9608
rect 4663 9605 4675 9639
rect 4617 9599 4675 9605
rect 5920 9577 5948 9676
rect 5994 9664 6000 9716
rect 6052 9664 6058 9716
rect 7466 9664 7472 9716
rect 7524 9664 7530 9716
rect 8202 9704 8208 9716
rect 8036 9676 8208 9704
rect 7484 9636 7512 9664
rect 8036 9645 8064 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9953 9707 10011 9713
rect 9953 9673 9965 9707
rect 9999 9704 10011 9707
rect 11514 9704 11520 9716
rect 9999 9676 11520 9704
rect 9999 9673 10011 9676
rect 9953 9667 10011 9673
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 11606 9664 11612 9716
rect 11664 9664 11670 9716
rect 8021 9639 8079 9645
rect 7484 9608 7788 9636
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4264 9540 4721 9568
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 2608 9364 2636 9463
rect 3234 9364 3240 9376
rect 2608 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4264 9364 4292 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7558 9568 7564 9580
rect 7515 9540 7564 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7760 9577 7788 9608
rect 8021 9605 8033 9639
rect 8067 9605 8079 9639
rect 8021 9599 8079 9605
rect 8478 9596 8484 9648
rect 8536 9596 8542 9648
rect 10502 9636 10508 9648
rect 9692 9608 10508 9636
rect 9692 9577 9720 9608
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 11146 9636 11152 9648
rect 10888 9608 11152 9636
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10686 9568 10692 9580
rect 10100 9540 10692 9568
rect 10100 9528 10106 9540
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 10888 9577 10916 9608
rect 11146 9596 11152 9608
rect 11204 9636 11210 9648
rect 12069 9639 12127 9645
rect 12069 9636 12081 9639
rect 11204 9608 12081 9636
rect 11204 9596 11210 9608
rect 12069 9605 12081 9608
rect 12115 9605 12127 9639
rect 12069 9599 12127 9605
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 10796 9500 10824 9531
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11422 9568 11428 9580
rect 11287 9540 11428 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11422 9528 11428 9540
rect 11480 9568 11486 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11480 9540 11805 9568
rect 11480 9528 11486 9540
rect 11793 9537 11805 9540
rect 11839 9568 11851 9571
rect 12710 9568 12716 9580
rect 11839 9540 12716 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 10980 9500 11008 9528
rect 10796 9472 11008 9500
rect 11885 9503 11943 9509
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9432 9551 9435
rect 10796 9432 10824 9472
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 9539 9404 10824 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10928 9404 10977 9432
rect 10928 9392 10934 9404
rect 10965 9401 10977 9404
rect 11011 9432 11023 9435
rect 11900 9432 11928 9463
rect 11011 9404 11928 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 3476 9336 4292 9364
rect 3476 9324 3482 9336
rect 4338 9324 4344 9376
rect 4396 9324 4402 9376
rect 7374 9324 7380 9376
rect 7432 9324 7438 9376
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10744 9336 11069 9364
rect 10744 9324 10750 9336
rect 11057 9333 11069 9336
rect 11103 9364 11115 9367
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11103 9336 12081 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 12069 9333 12081 9336
rect 12115 9364 12127 9367
rect 12618 9364 12624 9376
rect 12115 9336 12624 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 1104 9274 13340 9296
rect 1104 9222 2479 9274
rect 2531 9222 2543 9274
rect 2595 9222 2607 9274
rect 2659 9222 2671 9274
rect 2723 9222 2735 9274
rect 2787 9222 5538 9274
rect 5590 9222 5602 9274
rect 5654 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 8597 9274
rect 8649 9222 8661 9274
rect 8713 9222 8725 9274
rect 8777 9222 8789 9274
rect 8841 9222 8853 9274
rect 8905 9222 11656 9274
rect 11708 9222 11720 9274
rect 11772 9222 11784 9274
rect 11836 9222 11848 9274
rect 11900 9222 11912 9274
rect 11964 9222 13340 9274
rect 1104 9200 13340 9222
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 5506 9132 7205 9160
rect 4985 9095 5043 9101
rect 4985 9061 4997 9095
rect 5031 9092 5043 9095
rect 5031 9064 5212 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 5184 9036 5212 9064
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 5074 9024 5080 9036
rect 3292 8996 5080 9024
rect 3292 8984 3298 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5166 8984 5172 9036
rect 5224 8984 5230 9036
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 9024 5319 9027
rect 5506 9024 5534 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 7208 9092 7236 9123
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8297 9163 8355 9169
rect 7800 9132 8248 9160
rect 7800 9120 7806 9132
rect 7208 9064 7880 9092
rect 5307 8996 5534 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 3476 8928 3525 8956
rect 3476 8916 3482 8928
rect 3513 8925 3525 8928
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 4224 8959 4282 8965
rect 4224 8925 4236 8959
rect 4270 8956 4282 8959
rect 4338 8956 4344 8968
rect 4270 8928 4344 8956
rect 4270 8925 4282 8928
rect 4224 8919 4282 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5276 8956 5304 8987
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 7852 9033 7880 9064
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 6144 8996 7297 9024
rect 6144 8984 6150 8996
rect 7285 8993 7297 8996
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 7837 9027 7895 9033
rect 7837 8993 7849 9027
rect 7883 8993 7895 9027
rect 8220 9024 8248 9132
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8478 9160 8484 9172
rect 8343 9132 8484 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12342 9160 12348 9172
rect 12299 9132 12348 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 11514 9092 11520 9104
rect 11348 9064 11520 9092
rect 11348 9024 11376 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 8220 8996 11376 9024
rect 7837 8987 7895 8993
rect 4755 8928 5304 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 7374 8956 7380 8968
rect 6854 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 11348 8965 11376 8996
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7616 8928 8217 8956
rect 7616 8916 7622 8928
rect 8205 8925 8217 8928
rect 8251 8956 8263 8959
rect 11333 8959 11391 8965
rect 8251 8928 8340 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 2530 8860 2636 8888
rect 1486 8780 1492 8832
rect 1544 8780 1550 8832
rect 2608 8820 2636 8860
rect 2958 8848 2964 8900
rect 3016 8848 3022 8900
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4433 8891 4491 8897
rect 3844 8860 4384 8888
rect 3844 8848 3850 8860
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 2608 8792 3433 8820
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 4356 8829 4384 8860
rect 4433 8857 4445 8891
rect 4479 8888 4491 8891
rect 5166 8888 5172 8900
rect 4479 8860 5172 8888
rect 4479 8857 4491 8860
rect 4433 8851 4491 8857
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 5718 8848 5724 8900
rect 5776 8848 5782 8900
rect 8312 8832 8340 8928
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 12268 8956 12296 9123
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 11563 8928 12296 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3936 8792 4077 8820
rect 3936 8780 3942 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4065 8783 4123 8789
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4580 8792 4813 8820
rect 4580 8780 4586 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4801 8783 4859 8789
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 11422 8780 11428 8832
rect 11480 8780 11486 8832
rect 1104 8730 13499 8752
rect 1104 8678 4008 8730
rect 4060 8678 4072 8730
rect 4124 8678 4136 8730
rect 4188 8678 4200 8730
rect 4252 8678 4264 8730
rect 4316 8678 7067 8730
rect 7119 8678 7131 8730
rect 7183 8678 7195 8730
rect 7247 8678 7259 8730
rect 7311 8678 7323 8730
rect 7375 8678 10126 8730
rect 10178 8678 10190 8730
rect 10242 8678 10254 8730
rect 10306 8678 10318 8730
rect 10370 8678 10382 8730
rect 10434 8678 13185 8730
rect 13237 8678 13249 8730
rect 13301 8678 13313 8730
rect 13365 8678 13377 8730
rect 13429 8678 13441 8730
rect 13493 8678 13499 8730
rect 1104 8656 13499 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 2038 8616 2044 8628
rect 1544 8588 2044 8616
rect 1544 8576 1550 8588
rect 2038 8576 2044 8588
rect 2096 8616 2102 8628
rect 2096 8588 2774 8616
rect 2096 8576 2102 8588
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 2746 8548 2774 8588
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3016 8588 3249 8616
rect 3016 8576 3022 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3326 8576 3332 8628
rect 3384 8576 3390 8628
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 12342 8576 12348 8628
rect 12400 8576 12406 8628
rect 3513 8551 3571 8557
rect 2455 8520 2636 8548
rect 2746 8520 3004 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 2608 8489 2636 8520
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2317 8443 2375 8449
rect 2424 8452 2513 8480
rect 2332 8344 2360 8443
rect 2424 8424 2452 8452
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2774 8440 2780 8492
rect 2832 8440 2838 8492
rect 2866 8440 2872 8492
rect 2924 8440 2930 8492
rect 2976 8489 3004 8520
rect 3513 8517 3525 8551
rect 3559 8548 3571 8551
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3559 8520 3985 8548
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 4356 8548 4384 8576
rect 4614 8548 4620 8560
rect 3973 8511 4031 8517
rect 4172 8520 4620 8548
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3326 8480 3332 8492
rect 3007 8452 3332 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 4172 8489 4200 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 5224 8520 5534 8548
rect 5224 8508 5230 8520
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 5506 8480 5534 8520
rect 6362 8508 6368 8560
rect 6420 8508 6426 8560
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5506 8452 5917 8480
rect 4433 8443 4491 8449
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 8018 8480 8024 8492
rect 6227 8452 8024 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 2406 8372 2412 8424
rect 2464 8372 2470 8424
rect 3804 8412 3832 8440
rect 4448 8412 4476 8443
rect 2746 8384 4476 8412
rect 5920 8412 5948 8443
rect 8018 8440 8024 8452
rect 8076 8480 8082 8492
rect 8202 8480 8208 8492
rect 8076 8452 8208 8480
rect 8076 8440 8082 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12250 8480 12256 8492
rect 12115 8452 12256 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 10520 8412 10548 8440
rect 5920 8384 10548 8412
rect 2746 8344 2774 8384
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 2332 8316 2774 8344
rect 3878 8304 3884 8356
rect 3936 8304 3942 8356
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 2958 8276 2964 8288
rect 2832 8248 2964 8276
rect 2832 8236 2838 8248
rect 2958 8236 2964 8248
rect 3016 8276 3022 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 3016 8248 3525 8276
rect 3016 8236 3022 8248
rect 3513 8245 3525 8248
rect 3559 8245 3571 8279
rect 3513 8239 3571 8245
rect 7650 8236 7656 8288
rect 7708 8236 7714 8288
rect 12158 8236 12164 8288
rect 12216 8236 12222 8288
rect 1104 8186 13340 8208
rect 1104 8134 2479 8186
rect 2531 8134 2543 8186
rect 2595 8134 2607 8186
rect 2659 8134 2671 8186
rect 2723 8134 2735 8186
rect 2787 8134 5538 8186
rect 5590 8134 5602 8186
rect 5654 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 8597 8186
rect 8649 8134 8661 8186
rect 8713 8134 8725 8186
rect 8777 8134 8789 8186
rect 8841 8134 8853 8186
rect 8905 8134 11656 8186
rect 11708 8134 11720 8186
rect 11772 8134 11784 8186
rect 11836 8134 11848 8186
rect 11900 8134 11912 8186
rect 11964 8134 13340 8186
rect 1104 8112 13340 8134
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 2866 8072 2872 8084
rect 2639 8044 2872 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3786 8072 3792 8084
rect 3099 8044 3792 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5132 8044 5549 8072
rect 5132 8032 5138 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 12894 8032 12900 8084
rect 12952 8032 12958 8084
rect 2774 8004 2780 8016
rect 2240 7976 2780 8004
rect 2240 7945 2268 7976
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2884 7936 2912 8032
rect 2225 7899 2283 7905
rect 2516 7908 2912 7936
rect 2406 7828 2412 7880
rect 2464 7828 2470 7880
rect 2516 7877 2544 7908
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2961 7871 3019 7877
rect 2823 7840 2857 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3142 7868 3148 7880
rect 3007 7840 3148 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2792 7800 2820 7831
rect 3142 7828 3148 7840
rect 3200 7868 3206 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3200 7840 3249 7868
rect 3200 7828 3206 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6696 7840 7021 7868
rect 6696 7828 6702 7840
rect 7009 7837 7021 7840
rect 7055 7868 7067 7871
rect 7650 7868 7656 7880
rect 7055 7840 7656 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8478 7868 8484 7880
rect 8251 7840 8484 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 4356 7800 4384 7828
rect 2372 7772 4384 7800
rect 8128 7800 8156 7831
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9272 7840 9689 7868
rect 9272 7828 9278 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 8128 7772 8340 7800
rect 2372 7760 2378 7772
rect 8312 7744 8340 7772
rect 8938 7760 8944 7812
rect 8996 7760 9002 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9398 7800 9404 7812
rect 9171 7772 9404 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 12158 7760 12164 7812
rect 12216 7760 12222 7812
rect 2222 7692 2228 7744
rect 2280 7692 2286 7744
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 8294 7692 8300 7744
rect 8352 7692 8358 7744
rect 8386 7692 8392 7744
rect 8444 7692 8450 7744
rect 9306 7692 9312 7744
rect 9364 7692 9370 7744
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 1104 7642 13499 7664
rect 1104 7590 4008 7642
rect 4060 7590 4072 7642
rect 4124 7590 4136 7642
rect 4188 7590 4200 7642
rect 4252 7590 4264 7642
rect 4316 7590 7067 7642
rect 7119 7590 7131 7642
rect 7183 7590 7195 7642
rect 7247 7590 7259 7642
rect 7311 7590 7323 7642
rect 7375 7590 10126 7642
rect 10178 7590 10190 7642
rect 10242 7590 10254 7642
rect 10306 7590 10318 7642
rect 10370 7590 10382 7642
rect 10434 7590 13185 7642
rect 13237 7590 13249 7642
rect 13301 7590 13313 7642
rect 13365 7590 13377 7642
rect 13429 7590 13441 7642
rect 13493 7590 13499 7642
rect 1104 7568 13499 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2464 7500 2697 7528
rect 2464 7488 2470 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 2685 7491 2743 7497
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 6086 7460 6092 7472
rect 5767 7432 6092 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8404 7460 8432 7488
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 8404 7432 8769 7460
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 8757 7423 8815 7429
rect 9490 7420 9496 7472
rect 9548 7420 9554 7472
rect 11149 7463 11207 7469
rect 11149 7460 11161 7463
rect 10718 7432 11161 7460
rect 11149 7429 11161 7432
rect 11195 7429 11207 7463
rect 11149 7423 11207 7429
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2372 7364 2605 7392
rect 2372 7352 2378 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3142 7392 3148 7404
rect 2823 7364 3148 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 6181 7395 6239 7401
rect 6181 7392 6193 7395
rect 5920 7364 6193 7392
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 5920 7265 5948 7364
rect 6181 7361 6193 7364
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6564 7324 6592 7355
rect 9030 7352 9036 7404
rect 9088 7401 9094 7404
rect 9088 7395 9102 7401
rect 9090 7392 9102 7395
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 9090 7364 9229 7392
rect 9090 7361 9102 7364
rect 9088 7355 9102 7361
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11287 7364 12173 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 12161 7361 12173 7364
rect 12207 7392 12219 7395
rect 12207 7364 12296 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 9088 7352 9094 7355
rect 12268 7336 12296 7364
rect 6196 7296 6592 7324
rect 6196 7268 6224 7296
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 5040 7228 5365 7256
rect 5040 7216 5046 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7225 5963 7259
rect 5905 7219 5963 7225
rect 6178 7216 6184 7268
rect 6236 7216 6242 7268
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 4798 7188 4804 7200
rect 2832 7160 4804 7188
rect 2832 7148 2838 7160
rect 4798 7148 4804 7160
rect 4856 7188 4862 7200
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 4856 7160 5733 7188
rect 4856 7148 4862 7160
rect 5721 7157 5733 7160
rect 5767 7188 5779 7191
rect 5810 7188 5816 7200
rect 5767 7160 5816 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 5994 7148 6000 7200
rect 6052 7148 6058 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6604 7160 6653 7188
rect 6604 7148 6610 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7558 7188 7564 7200
rect 7331 7160 7564 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 10134 7188 10140 7200
rect 9548 7160 10140 7188
rect 9548 7148 9554 7160
rect 10134 7148 10140 7160
rect 10192 7188 10198 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10192 7160 10977 7188
rect 10192 7148 10198 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12253 7191 12311 7197
rect 12253 7188 12265 7191
rect 12216 7160 12265 7188
rect 12216 7148 12222 7160
rect 12253 7157 12265 7160
rect 12299 7157 12311 7191
rect 12253 7151 12311 7157
rect 1104 7098 13340 7120
rect 1104 7046 2479 7098
rect 2531 7046 2543 7098
rect 2595 7046 2607 7098
rect 2659 7046 2671 7098
rect 2723 7046 2735 7098
rect 2787 7046 5538 7098
rect 5590 7046 5602 7098
rect 5654 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 8597 7098
rect 8649 7046 8661 7098
rect 8713 7046 8725 7098
rect 8777 7046 8789 7098
rect 8841 7046 8853 7098
rect 8905 7046 11656 7098
rect 11708 7046 11720 7098
rect 11772 7046 11784 7098
rect 11836 7046 11848 7098
rect 11900 7046 11912 7098
rect 11964 7046 13340 7098
rect 1104 7024 13340 7046
rect 1660 6987 1718 6993
rect 1660 6953 1672 6987
rect 1706 6984 1718 6987
rect 2222 6984 2228 6996
rect 1706 6956 2228 6984
rect 1706 6953 1718 6956
rect 1660 6947 1718 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 5960 6956 8401 6984
rect 5960 6944 5966 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 1394 6808 1400 6860
rect 1452 6808 1458 6860
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5500 6820 5549 6848
rect 5500 6808 5506 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5902 6848 5908 6860
rect 5859 6820 5908 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 8404 6848 8432 6947
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 8536 6956 8585 6984
rect 8536 6944 8542 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 8573 6947 8631 6953
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9214 6984 9220 6996
rect 9171 6956 9220 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6953 9367 6987
rect 9309 6947 9367 6953
rect 9324 6916 9352 6947
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9953 6987 10011 6993
rect 9953 6984 9965 6987
rect 9640 6956 9965 6984
rect 9640 6944 9646 6956
rect 9953 6953 9965 6956
rect 9999 6953 10011 6987
rect 9953 6947 10011 6953
rect 10597 6987 10655 6993
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 10778 6984 10784 6996
rect 10643 6956 10784 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 10612 6916 10640 6947
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 9048 6888 10640 6916
rect 9048 6848 9076 6888
rect 11146 6848 11152 6860
rect 8404 6820 9076 6848
rect 9324 6820 11152 6848
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3418 6780 3424 6792
rect 3016 6752 3424 6780
rect 3016 6740 3022 6752
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7668 6752 7757 6780
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 2898 6684 3341 6712
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3752 6684 4169 6712
rect 3752 6672 3758 6684
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4157 6675 4215 6681
rect 4338 6672 4344 6724
rect 4396 6672 4402 6724
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5077 6715 5135 6721
rect 5077 6712 5089 6715
rect 4488 6684 5089 6712
rect 4488 6672 4494 6684
rect 5077 6681 5089 6684
rect 5123 6681 5135 6715
rect 5077 6675 5135 6681
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5350 6712 5356 6724
rect 5307 6684 5356 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 6086 6712 6092 6724
rect 5491 6684 6092 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 6546 6672 6552 6724
rect 6604 6672 6610 6724
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 4522 6604 4528 6656
rect 4580 6604 4586 6656
rect 4706 6604 4712 6656
rect 4764 6604 4770 6656
rect 5368 6644 5396 6672
rect 7668 6656 7696 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7975 6752 8033 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8021 6749 8033 6752
rect 8067 6780 8079 6783
rect 8938 6780 8944 6792
rect 8067 6752 8944 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9324 6780 9352 6820
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 9088 6752 9352 6780
rect 9677 6783 9735 6789
rect 9088 6740 9094 6752
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 9766 6780 9772 6792
rect 9723 6752 9772 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 9916 6752 10241 6780
rect 9916 6740 9922 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10229 6743 10287 6749
rect 10796 6752 10885 6780
rect 9306 6672 9312 6724
rect 9364 6672 9370 6724
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 5368 6616 7297 6644
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 9784 6653 9812 6740
rect 10134 6672 10140 6724
rect 10192 6672 10198 6724
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 9927 6647 9985 6653
rect 9927 6613 9939 6647
rect 9973 6644 9985 6647
rect 10042 6644 10048 6656
rect 9973 6616 10048 6644
rect 9973 6613 9985 6616
rect 9927 6607 9985 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 10594 6604 10600 6656
rect 10652 6604 10658 6656
rect 10796 6653 10824 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11425 6715 11483 6721
rect 11425 6712 11437 6715
rect 11072 6684 11437 6712
rect 11072 6653 11100 6684
rect 11425 6681 11437 6684
rect 11471 6681 11483 6715
rect 11425 6675 11483 6681
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 12894 6604 12900 6656
rect 12952 6604 12958 6656
rect 1104 6554 13499 6576
rect 1104 6502 4008 6554
rect 4060 6502 4072 6554
rect 4124 6502 4136 6554
rect 4188 6502 4200 6554
rect 4252 6502 4264 6554
rect 4316 6502 7067 6554
rect 7119 6502 7131 6554
rect 7183 6502 7195 6554
rect 7247 6502 7259 6554
rect 7311 6502 7323 6554
rect 7375 6502 10126 6554
rect 10178 6502 10190 6554
rect 10242 6502 10254 6554
rect 10306 6502 10318 6554
rect 10370 6502 10382 6554
rect 10434 6502 13185 6554
rect 13237 6502 13249 6554
rect 13301 6502 13313 6554
rect 13365 6502 13377 6554
rect 13429 6502 13441 6554
rect 13493 6502 13499 6554
rect 1104 6480 13499 6502
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4430 6440 4436 6452
rect 3927 6412 4436 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 7650 6440 7656 6452
rect 5040 6412 7656 6440
rect 5040 6400 5046 6412
rect 7650 6400 7656 6412
rect 7708 6440 7714 6452
rect 7708 6412 8248 6440
rect 7708 6400 7714 6412
rect 4033 6375 4091 6381
rect 4033 6372 4045 6375
rect 3896 6344 4045 6372
rect 3896 6316 3924 6344
rect 4033 6341 4045 6344
rect 4079 6341 4091 6375
rect 4249 6375 4307 6381
rect 4249 6372 4261 6375
rect 4033 6335 4091 6341
rect 4172 6344 4261 6372
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 2869 6307 2927 6313
rect 2639 6276 2774 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2746 6236 2774 6276
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 2958 6304 2964 6316
rect 2915 6276 2964 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6304 3571 6307
rect 3878 6304 3884 6316
rect 3559 6276 3884 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 3050 6236 3056 6248
rect 2746 6208 3056 6236
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3375 6208 3832 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3804 6112 3832 6208
rect 4172 6168 4200 6344
rect 4249 6341 4261 6344
rect 4295 6372 4307 6375
rect 4338 6372 4344 6384
rect 4295 6344 4344 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 4724 6372 4752 6400
rect 5902 6372 5908 6384
rect 4663 6344 4752 6372
rect 5842 6344 5908 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 7558 6332 7564 6384
rect 7616 6332 7622 6384
rect 8220 6381 8248 6412
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8444 6412 8585 6440
rect 8444 6400 8450 6412
rect 8573 6409 8585 6412
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 9490 6400 9496 6452
rect 9548 6400 9554 6452
rect 9766 6400 9772 6452
rect 9824 6400 9830 6452
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10594 6440 10600 6452
rect 10367 6412 10600 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 8205 6375 8263 6381
rect 8205 6341 8217 6375
rect 8251 6372 8263 6375
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 8251 6344 9689 6372
rect 8251 6341 8263 6344
rect 8205 6335 8263 6341
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 9784 6372 9812 6400
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 9784 6344 9965 6372
rect 9677 6335 9735 6341
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 10137 6375 10195 6381
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 12894 6372 12900 6384
rect 10183 6344 12900 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 7576 6304 7604 6332
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 7576 6276 8401 6304
rect 8389 6273 8401 6276
rect 8435 6304 8447 6307
rect 9582 6304 9588 6316
rect 8435 6276 9588 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9692 6304 9720 6335
rect 10042 6304 10048 6316
rect 9692 6276 10048 6304
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 4338 6236 4344 6248
rect 4396 6245 4402 6248
rect 4306 6208 4344 6236
rect 4338 6196 4344 6208
rect 4396 6199 4406 6245
rect 5258 6236 5264 6248
rect 4448 6208 5264 6236
rect 4396 6196 4402 6199
rect 4448 6168 4476 6208
rect 5258 6196 5264 6208
rect 5316 6236 5322 6248
rect 6089 6239 6147 6245
rect 6089 6236 6101 6239
rect 5316 6208 6101 6236
rect 5316 6196 5322 6208
rect 6089 6205 6101 6208
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9766 6236 9772 6248
rect 9355 6208 9772 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9766 6196 9772 6208
rect 9824 6236 9830 6248
rect 10152 6236 10180 6335
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 9824 6208 10180 6236
rect 9824 6196 9830 6208
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 4172 6140 4476 6168
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2188 6072 2421 6100
rect 2188 6060 2194 6072
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3694 6100 3700 6112
rect 3384 6072 3700 6100
rect 3384 6060 3390 6072
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3844 6072 4077 6100
rect 3844 6060 3850 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4798 6100 4804 6112
rect 4396 6072 4804 6100
rect 4396 6060 4402 6072
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 8294 6100 8300 6112
rect 6236 6072 8300 6100
rect 6236 6060 6242 6072
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 1104 6010 13340 6032
rect 1104 5958 2479 6010
rect 2531 5958 2543 6010
rect 2595 5958 2607 6010
rect 2659 5958 2671 6010
rect 2723 5958 2735 6010
rect 2787 5958 5538 6010
rect 5590 5958 5602 6010
rect 5654 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 8597 6010
rect 8649 5958 8661 6010
rect 8713 5958 8725 6010
rect 8777 5958 8789 6010
rect 8841 5958 8853 6010
rect 8905 5958 11656 6010
rect 11708 5958 11720 6010
rect 11772 5958 11784 6010
rect 11836 5958 11848 6010
rect 11900 5958 11912 6010
rect 11964 5958 13340 6010
rect 1104 5936 13340 5958
rect 4246 5896 4252 5908
rect 1504 5868 4252 5896
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1504 5769 1532 5868
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4890 5896 4896 5908
rect 4571 5868 4896 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 6328 5868 6469 5896
rect 6328 5856 6334 5868
rect 6457 5865 6469 5868
rect 6503 5896 6515 5899
rect 7466 5896 7472 5908
rect 6503 5868 7472 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 7947 5899 8005 5905
rect 7947 5865 7959 5899
rect 7993 5896 8005 5899
rect 8754 5896 8760 5908
rect 7993 5868 8760 5896
rect 7993 5865 8005 5868
rect 7947 5859 8005 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 4264 5828 4292 5856
rect 5442 5828 5448 5840
rect 4264 5800 5448 5828
rect 1489 5763 1547 5769
rect 1489 5760 1501 5763
rect 1452 5732 1501 5760
rect 1452 5720 1458 5732
rect 1489 5729 1501 5732
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2130 5760 2136 5772
rect 1811 5732 2136 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5760 4031 5763
rect 4430 5760 4436 5772
rect 4019 5732 4436 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4522 5720 4528 5772
rect 4580 5720 4586 5772
rect 4632 5769 4660 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 5460 5760 5488 5788
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 5460 5732 8217 5760
rect 4617 5723 4675 5729
rect 8205 5729 8217 5732
rect 8251 5760 8263 5763
rect 9030 5760 9036 5772
rect 8251 5732 9036 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4540 5624 4568 5720
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6638 5692 6644 5704
rect 6411 5664 6644 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8389 5627 8447 5633
rect 4387 5596 4568 5624
rect 7498 5596 7604 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3694 5556 3700 5568
rect 3283 5528 3700 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 7576 5556 7604 5596
rect 8389 5593 8401 5627
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 8404 5556 8432 5587
rect 7576 5528 8432 5556
rect 1104 5466 13499 5488
rect 1104 5414 4008 5466
rect 4060 5414 4072 5466
rect 4124 5414 4136 5466
rect 4188 5414 4200 5466
rect 4252 5414 4264 5466
rect 4316 5414 7067 5466
rect 7119 5414 7131 5466
rect 7183 5414 7195 5466
rect 7247 5414 7259 5466
rect 7311 5414 7323 5466
rect 7375 5414 10126 5466
rect 10178 5414 10190 5466
rect 10242 5414 10254 5466
rect 10306 5414 10318 5466
rect 10370 5414 10382 5466
rect 10434 5414 13185 5466
rect 13237 5414 13249 5466
rect 13301 5414 13313 5466
rect 13365 5414 13377 5466
rect 13429 5414 13441 5466
rect 13493 5414 13499 5466
rect 1104 5392 13499 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 3050 5352 3056 5364
rect 2823 5324 3056 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 4982 5312 4988 5364
rect 5040 5312 5046 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5316 5324 5365 5352
rect 5316 5312 5322 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5902 5352 5908 5364
rect 5767 5324 5908 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 9490 5312 9496 5364
rect 9548 5312 9554 5364
rect 9766 5312 9772 5364
rect 9824 5312 9830 5364
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 11165 5355 11223 5361
rect 11165 5352 11177 5355
rect 10796 5324 11177 5352
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 3007 5256 3801 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3789 5253 3801 5256
rect 3835 5253 3847 5287
rect 3789 5247 3847 5253
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 4157 5287 4215 5293
rect 4157 5284 4169 5287
rect 3936 5256 4169 5284
rect 3936 5244 3942 5256
rect 4157 5253 4169 5256
rect 4203 5284 4215 5287
rect 5169 5287 5227 5293
rect 5169 5284 5181 5287
rect 4203 5256 5181 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 5169 5253 5181 5256
rect 5215 5253 5227 5287
rect 5169 5247 5227 5253
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6914 5284 6920 5296
rect 5592 5256 6920 5284
rect 5592 5244 5598 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 8294 5293 8300 5296
rect 8271 5287 8300 5293
rect 8271 5253 8283 5287
rect 8271 5247 8300 5253
rect 8294 5244 8300 5247
rect 8352 5244 8358 5296
rect 8389 5287 8447 5293
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 9122 5284 9128 5296
rect 8435 5256 9128 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2148 5024 2176 5179
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3752 5188 3985 5216
rect 3752 5176 3758 5188
rect 3973 5185 3985 5188
rect 4019 5216 4031 5219
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4019 5188 5273 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6086 5216 6092 5228
rect 5859 5188 6092 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2958 5148 2964 5160
rect 2455 5120 2964 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2958 5108 2964 5120
rect 3016 5148 3022 5160
rect 5828 5148 5856 5179
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 9214 5216 9220 5228
rect 8619 5188 9220 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9508 5216 9536 5312
rect 9784 5225 9812 5312
rect 9355 5188 9536 5216
rect 9769 5219 9827 5225
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 9769 5185 9781 5219
rect 9815 5185 9827 5219
rect 9876 5216 9904 5312
rect 10505 5287 10563 5293
rect 10505 5284 10517 5287
rect 10244 5256 10517 5284
rect 10244 5225 10272 5256
rect 10505 5253 10517 5256
rect 10551 5253 10563 5287
rect 10505 5247 10563 5253
rect 10796 5228 10824 5324
rect 11165 5321 11177 5324
rect 11211 5321 11223 5355
rect 11165 5315 11223 5321
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 10965 5287 11023 5293
rect 10965 5253 10977 5287
rect 11011 5284 11023 5287
rect 11011 5256 11284 5284
rect 11011 5253 11023 5256
rect 10965 5247 11023 5253
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9876 5188 10241 5216
rect 9769 5179 9827 5185
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 10686 5216 10692 5228
rect 10459 5188 10692 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 11256 5160 11284 5256
rect 11348 5216 11376 5315
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11348 5188 11713 5216
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 3016 5120 5856 5148
rect 8021 5151 8079 5157
rect 3016 5108 3022 5120
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 8067 5120 8125 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 11238 5148 11244 5160
rect 10367 5120 11244 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 12176 5148 12204 5176
rect 12434 5148 12440 5160
rect 12176 5120 12440 5148
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 12176 5080 12204 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 5224 5052 12204 5080
rect 5224 5040 5230 5052
rect 2130 4972 2136 5024
rect 2188 4972 2194 5024
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 4338 5012 4344 5024
rect 3007 4984 4344 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 9217 5015 9275 5021
rect 9217 4981 9229 5015
rect 9263 5012 9275 5015
rect 9398 5012 9404 5024
rect 9263 4984 9404 5012
rect 9263 4981 9275 4984
rect 9217 4975 9275 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 9766 5012 9772 5024
rect 9723 4984 9772 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10873 5015 10931 5021
rect 10873 4981 10885 5015
rect 10919 5012 10931 5015
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10919 4984 11161 5012
rect 10919 4981 10931 4984
rect 10873 4975 10931 4981
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 12216 4984 12265 5012
rect 12216 4972 12222 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 1104 4922 13340 4944
rect 1104 4870 2479 4922
rect 2531 4870 2543 4922
rect 2595 4870 2607 4922
rect 2659 4870 2671 4922
rect 2723 4870 2735 4922
rect 2787 4870 5538 4922
rect 5590 4870 5602 4922
rect 5654 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 8597 4922
rect 8649 4870 8661 4922
rect 8713 4870 8725 4922
rect 8777 4870 8789 4922
rect 8841 4870 8853 4922
rect 8905 4870 11656 4922
rect 11708 4870 11720 4922
rect 11772 4870 11784 4922
rect 11836 4870 11848 4922
rect 11900 4870 11912 4922
rect 11964 4870 13340 4922
rect 1104 4848 13340 4870
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 9272 4780 10701 4808
rect 9272 4768 9278 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 5166 4672 5172 4684
rect 3007 4644 5172 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11514 4672 11520 4684
rect 11471 4644 11520 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 2130 4604 2136 4616
rect 1397 4567 1455 4573
rect 1596 4576 2136 4604
rect 1596 4477 1624 4576
rect 2130 4564 2136 4576
rect 2188 4604 2194 4616
rect 2685 4607 2743 4613
rect 2685 4604 2697 4607
rect 2188 4576 2697 4604
rect 2188 4564 2194 4576
rect 2685 4573 2697 4576
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 10919 4576 11100 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 10704 4536 10732 4564
rect 10962 4536 10968 4548
rect 10704 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11072 4480 11100 4576
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 12158 4496 12164 4548
rect 12216 4496 12222 4548
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 11054 4428 11060 4480
rect 11112 4428 11118 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 11388 4440 12909 4468
rect 11388 4428 11394 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 1104 4378 13499 4400
rect 1104 4326 4008 4378
rect 4060 4326 4072 4378
rect 4124 4326 4136 4378
rect 4188 4326 4200 4378
rect 4252 4326 4264 4378
rect 4316 4326 7067 4378
rect 7119 4326 7131 4378
rect 7183 4326 7195 4378
rect 7247 4326 7259 4378
rect 7311 4326 7323 4378
rect 7375 4326 10126 4378
rect 10178 4326 10190 4378
rect 10242 4326 10254 4378
rect 10306 4326 10318 4378
rect 10370 4326 10382 4378
rect 10434 4326 13185 4378
rect 13237 4326 13249 4378
rect 13301 4326 13313 4378
rect 13365 4326 13377 4378
rect 13429 4326 13441 4378
rect 13493 4326 13499 4378
rect 1104 4304 13499 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 7650 4264 7656 4276
rect 3660 4236 6224 4264
rect 3660 4224 3666 4236
rect 2792 4168 3004 4196
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4126 2283 4131
rect 2314 4126 2320 4140
rect 2271 4098 2320 4126
rect 2271 4097 2283 4098
rect 2225 4091 2283 4097
rect 2314 4088 2320 4098
rect 2372 4128 2378 4140
rect 2792 4128 2820 4168
rect 2372 4100 2820 4128
rect 2372 4088 2378 4100
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 2976 4128 3004 4168
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 5629 4199 5687 4205
rect 4120 4168 5028 4196
rect 4120 4156 4126 4168
rect 4540 4137 4568 4168
rect 5000 4140 5028 4168
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5675 4168 5856 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 4525 4131 4583 4137
rect 2976 4100 4476 4128
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 2096 4032 3556 4060
rect 2096 4020 2102 4032
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3992 2651 3995
rect 3142 3992 3148 4004
rect 2639 3964 3148 3992
rect 2639 3961 2651 3964
rect 2593 3955 2651 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3528 3992 3556 4032
rect 3694 4020 3700 4072
rect 3752 4020 3758 4072
rect 4448 4060 4476 4100
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5123 4100 5733 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5828 4128 5856 4168
rect 6086 4128 6092 4140
rect 5828 4100 6092 4128
rect 5721 4091 5779 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6196 4128 6224 4236
rect 7208 4236 7656 4264
rect 7208 4137 7236 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8536 4236 8585 4264
rect 8536 4224 8542 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 10229 4267 10287 4273
rect 10229 4233 10241 4267
rect 10275 4264 10287 4267
rect 10778 4264 10784 4276
rect 10275 4236 10784 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11330 4264 11336 4276
rect 11020 4236 11336 4264
rect 11020 4224 11026 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 7484 4168 8524 4196
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6196 4100 6929 4128
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7340 4100 7389 4128
rect 7340 4088 7346 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 5813 4063 5871 4069
rect 3804 4032 4292 4060
rect 4448 4032 5396 4060
rect 3804 3992 3832 4032
rect 4264 4004 4292 4032
rect 3252 3964 3464 3992
rect 3528 3964 3832 3992
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2866 3924 2872 3936
rect 2731 3896 2872 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 2958 3884 2964 3936
rect 3016 3884 3022 3936
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3252 3924 3280 3964
rect 3108 3896 3280 3924
rect 3108 3884 3114 3896
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 3436 3924 3464 3964
rect 4062 3952 4068 4004
rect 4120 3952 4126 4004
rect 4246 3952 4252 4004
rect 4304 3952 4310 4004
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 4764 3964 5212 3992
rect 4764 3952 4770 3964
rect 3694 3924 3700 3936
rect 3436 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4080 3924 4108 3952
rect 3844 3896 4108 3924
rect 4157 3927 4215 3933
rect 3844 3884 3850 3896
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4338 3924 4344 3936
rect 4203 3896 4344 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 5074 3924 5080 3936
rect 4663 3896 5080 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5184 3933 5212 3964
rect 5258 3952 5264 4004
rect 5316 3952 5322 4004
rect 5368 3992 5396 4032
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5902 4060 5908 4072
rect 5859 4032 5908 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 5994 4020 6000 4072
rect 6052 4020 6058 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6696 4032 6745 4060
rect 6696 4020 6702 4032
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7484 4060 7512 4168
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 6880 4032 7512 4060
rect 6880 4020 6886 4032
rect 7009 3995 7067 4001
rect 7009 3992 7021 3995
rect 5368 3964 7021 3992
rect 7009 3961 7021 3964
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 7098 3952 7104 4004
rect 7156 3952 7162 4004
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6638 3924 6644 3936
rect 5951 3896 6644 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 7576 3924 7604 4091
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 8168 4100 8217 4128
rect 8168 4088 8174 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8312 4060 8340 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8496 4128 8524 4168
rect 8772 4168 8984 4196
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8496 4100 8677 4128
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8772 4060 8800 4168
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8312 4032 8800 4060
rect 7650 3952 7656 4004
rect 7708 3952 7714 4004
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8864 3992 8892 4091
rect 8956 4060 8984 4168
rect 9122 4156 9128 4208
rect 9180 4196 9186 4208
rect 9180 4168 9904 4196
rect 9180 4156 9186 4168
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9088 4100 9413 4128
rect 9088 4088 9094 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 9876 4128 9904 4168
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11149 4199 11207 4205
rect 11149 4196 11161 4199
rect 11112 4168 11161 4196
rect 11112 4156 11118 4168
rect 11149 4165 11161 4168
rect 11195 4196 11207 4199
rect 11195 4168 12940 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 12912 4140 12940 4168
rect 10379 4131 10437 4137
rect 10379 4128 10391 4131
rect 9876 4100 10391 4128
rect 10379 4097 10391 4100
rect 10425 4128 10437 4131
rect 10425 4100 10548 4128
rect 10425 4097 10437 4100
rect 10379 4091 10437 4097
rect 9784 4060 9812 4088
rect 8956 4032 9812 4060
rect 10520 4004 10548 4100
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 11747 4100 12357 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12894 4088 12900 4140
rect 12952 4088 12958 4140
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 7975 3964 8892 3992
rect 9048 3964 10364 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 6788 3896 7604 3924
rect 7668 3924 7696 3952
rect 9048 3936 9076 3964
rect 8754 3924 8760 3936
rect 7668 3896 8760 3924
rect 6788 3884 6794 3896
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 8938 3924 8944 3936
rect 8895 3896 8944 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9030 3884 9036 3936
rect 9088 3884 9094 3936
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 10336 3924 10364 3964
rect 10502 3952 10508 4004
rect 10560 3952 10566 4004
rect 10796 3992 10824 4023
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11296 4032 11621 4060
rect 11296 4020 11302 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 10796 3964 11161 3992
rect 11149 3961 11161 3964
rect 11195 3961 11207 3995
rect 11149 3955 11207 3961
rect 10778 3924 10784 3936
rect 10336 3896 10784 3924
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 12066 3884 12072 3936
rect 12124 3884 12130 3936
rect 1104 3834 13340 3856
rect 1104 3782 2479 3834
rect 2531 3782 2543 3834
rect 2595 3782 2607 3834
rect 2659 3782 2671 3834
rect 2723 3782 2735 3834
rect 2787 3782 5538 3834
rect 5590 3782 5602 3834
rect 5654 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 8597 3834
rect 8649 3782 8661 3834
rect 8713 3782 8725 3834
rect 8777 3782 8789 3834
rect 8841 3782 8853 3834
rect 8905 3782 11656 3834
rect 11708 3782 11720 3834
rect 11772 3782 11784 3834
rect 11836 3782 11848 3834
rect 11900 3782 11912 3834
rect 11964 3782 13340 3834
rect 1104 3760 13340 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1719 3692 2329 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 2317 3683 2375 3689
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3720 2743 3723
rect 2866 3720 2872 3732
rect 2731 3692 2872 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3652 2007 3655
rect 2222 3652 2228 3664
rect 1995 3624 2228 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 1578 3584 1584 3596
rect 1412 3556 1584 3584
rect 1412 3525 1440 3556
rect 1578 3544 1584 3556
rect 1636 3584 1642 3596
rect 1964 3584 1992 3615
rect 2222 3612 2228 3624
rect 2280 3612 2286 3664
rect 1636 3556 1992 3584
rect 1636 3544 1642 3556
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 2332 3584 2360 3683
rect 2866 3680 2872 3692
rect 2924 3720 2930 3732
rect 4525 3723 4583 3729
rect 2924 3692 4200 3720
rect 2924 3680 2930 3692
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3652 2559 3655
rect 2547 3624 3280 3652
rect 2547 3621 2559 3624
rect 2501 3615 2559 3621
rect 3142 3584 3148 3596
rect 2332 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3485 1455 3519
rect 2056 3516 2084 3544
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2056 3488 2605 3516
rect 1397 3479 1455 3485
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 2961 3451 3019 3457
rect 2961 3448 2973 3451
rect 1872 3420 2973 3448
rect 1872 3389 1900 3420
rect 2961 3417 2973 3420
rect 3007 3417 3019 3451
rect 3252 3448 3280 3624
rect 3326 3612 3332 3664
rect 3384 3612 3390 3664
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3878 3652 3884 3664
rect 3559 3624 3884 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 3878 3612 3884 3624
rect 3936 3652 3942 3664
rect 3936 3624 4108 3652
rect 3936 3612 3942 3624
rect 3344 3584 3372 3612
rect 4080 3593 4108 3624
rect 4172 3593 4200 3692
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 4798 3720 4804 3732
rect 4571 3692 4804 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 6822 3720 6828 3732
rect 5583 3692 6828 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7006 3680 7012 3732
rect 7064 3680 7070 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7156 3692 7389 3720
rect 7156 3680 7162 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8076 3692 8953 3720
rect 8076 3680 8082 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 9306 3720 9312 3732
rect 8941 3683 8999 3689
rect 9048 3692 9312 3720
rect 5092 3652 5120 3680
rect 5442 3652 5448 3664
rect 5092 3624 5448 3652
rect 4065 3587 4123 3593
rect 3344 3556 3832 3584
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3602 3516 3608 3528
rect 3467 3488 3608 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 3804 3525 3832 3556
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 5092 3584 5120 3624
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 5721 3655 5779 3661
rect 5721 3652 5733 3655
rect 5500 3624 5733 3652
rect 5500 3612 5506 3624
rect 5721 3621 5733 3624
rect 5767 3621 5779 3655
rect 6086 3652 6092 3664
rect 5721 3615 5779 3621
rect 5828 3624 6092 3652
rect 4157 3547 4215 3553
rect 4448 3556 5028 3584
rect 5092 3556 5212 3584
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 3988 3448 4016 3479
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 4304 3488 4353 3516
rect 4304 3476 4310 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 3252 3420 4016 3448
rect 2961 3411 3019 3417
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 2096 3352 2329 3380
rect 2096 3340 2102 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2866 3340 2872 3392
rect 2924 3340 2930 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 4448 3380 4476 3556
rect 5000 3525 5028 3556
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 3375 3352 4476 3380
rect 4816 3380 4844 3479
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5184 3525 5212 3556
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5828 3525 5856 3624
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 6365 3655 6423 3661
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 7742 3652 7748 3664
rect 6411 3624 7748 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 7834 3612 7840 3664
rect 7892 3652 7898 3664
rect 9048 3652 9076 3692
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9401 3723 9459 3729
rect 9401 3689 9413 3723
rect 9447 3720 9459 3723
rect 10042 3720 10048 3732
rect 9447 3692 10048 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10229 3723 10287 3729
rect 10229 3689 10241 3723
rect 10275 3720 10287 3723
rect 10686 3720 10692 3732
rect 10275 3692 10692 3720
rect 10275 3689 10287 3692
rect 10229 3683 10287 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10928 3692 10977 3720
rect 10928 3680 10934 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 10965 3683 11023 3689
rect 12894 3680 12900 3732
rect 12952 3680 12958 3732
rect 9766 3652 9772 3664
rect 7892 3624 8156 3652
rect 7892 3612 7898 3624
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3584 5963 3587
rect 5994 3584 6000 3596
rect 5951 3556 6000 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6270 3584 6276 3596
rect 6104 3556 6276 3584
rect 6104 3525 6132 3556
rect 6270 3544 6276 3556
rect 6328 3584 6334 3596
rect 6730 3584 6736 3596
rect 6328 3556 6736 3584
rect 6328 3544 6334 3556
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6914 3544 6920 3596
rect 6972 3544 6978 3596
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 7208 3556 7972 3584
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 5368 3448 5396 3479
rect 6196 3448 6224 3479
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6420 3488 6469 3516
rect 6420 3476 6426 3488
rect 6457 3485 6469 3488
rect 6503 3516 6515 3519
rect 6932 3516 6960 3544
rect 7208 3525 7236 3556
rect 6503 3488 6960 3516
rect 7193 3519 7251 3525
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7594 3519 7652 3525
rect 7594 3516 7606 3519
rect 7340 3488 7606 3516
rect 7340 3476 7346 3488
rect 7594 3485 7606 3488
rect 7640 3485 7652 3519
rect 7944 3516 7972 3556
rect 8018 3544 8024 3596
rect 8076 3544 8082 3596
rect 8128 3593 8156 3624
rect 8772 3624 9076 3652
rect 9232 3624 9772 3652
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8772 3584 8800 3624
rect 8720 3556 8800 3584
rect 8720 3544 8726 3556
rect 8772 3525 8800 3556
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 9030 3544 9036 3596
rect 9088 3544 9094 3596
rect 8389 3519 8447 3525
rect 7944 3488 8156 3516
rect 7594 3479 7652 3485
rect 5368 3420 6224 3448
rect 6914 3408 6920 3460
rect 6972 3408 6978 3460
rect 8128 3448 8156 3488
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8757 3519 8815 3525
rect 8435 3488 8708 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8404 3448 8432 3479
rect 8128 3420 8432 3448
rect 8481 3451 8539 3457
rect 8481 3417 8493 3451
rect 8527 3417 8539 3451
rect 8481 3411 8539 3417
rect 5534 3380 5540 3392
rect 4816 3352 5540 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 7742 3380 7748 3392
rect 7699 3352 7748 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8202 3340 8208 3392
rect 8260 3340 8266 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8500 3380 8528 3411
rect 8570 3408 8576 3460
rect 8628 3408 8634 3460
rect 8680 3448 8708 3488
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8846 3448 8852 3460
rect 8680 3420 8852 3448
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 8956 3448 8984 3544
rect 9048 3516 9076 3544
rect 9232 3528 9260 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 9600 3556 10517 3584
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9048 3488 9137 3516
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9214 3476 9220 3528
rect 9272 3476 9278 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9600 3525 9628 3556
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10888 3584 10916 3680
rect 10505 3547 10563 3553
rect 10612 3556 10916 3584
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9824 3488 9965 3516
rect 9824 3476 9830 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10042 3476 10048 3528
rect 10100 3525 10106 3528
rect 10612 3525 10640 3556
rect 11146 3544 11152 3596
rect 11204 3544 11210 3596
rect 10100 3516 10108 3525
rect 10413 3519 10471 3525
rect 10100 3488 10145 3516
rect 10100 3479 10108 3488
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10100 3476 10106 3479
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 8956 3420 9873 3448
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 10428 3448 10456 3479
rect 10870 3476 10876 3528
rect 10928 3476 10934 3528
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 12526 3476 12532 3528
rect 12584 3476 12590 3528
rect 10980 3448 11008 3476
rect 10428 3420 11008 3448
rect 11425 3451 11483 3457
rect 9861 3411 9919 3417
rect 11425 3417 11437 3451
rect 11471 3417 11483 3451
rect 11425 3411 11483 3417
rect 9398 3380 9404 3392
rect 8352 3352 9404 3380
rect 8352 3340 8358 3352
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 11440 3380 11468 3411
rect 12158 3380 12164 3392
rect 11440 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 1104 3290 13499 3312
rect 1104 3238 4008 3290
rect 4060 3238 4072 3290
rect 4124 3238 4136 3290
rect 4188 3238 4200 3290
rect 4252 3238 4264 3290
rect 4316 3238 7067 3290
rect 7119 3238 7131 3290
rect 7183 3238 7195 3290
rect 7247 3238 7259 3290
rect 7311 3238 7323 3290
rect 7375 3238 10126 3290
rect 10178 3238 10190 3290
rect 10242 3238 10254 3290
rect 10306 3238 10318 3290
rect 10370 3238 10382 3290
rect 10434 3238 13185 3290
rect 13237 3238 13249 3290
rect 13301 3238 13313 3290
rect 13365 3238 13377 3290
rect 13429 3238 13441 3290
rect 13493 3238 13499 3290
rect 1104 3216 13499 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2924 3148 2973 3176
rect 2924 3136 2930 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3050 3136 3056 3188
rect 3108 3136 3114 3188
rect 4246 3176 4252 3188
rect 3252 3148 4252 3176
rect 3252 3108 3280 3148
rect 4080 3117 4108 3148
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4338 3136 4344 3188
rect 4396 3136 4402 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4890 3176 4896 3188
rect 4479 3148 4896 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5442 3136 5448 3188
rect 5500 3136 5506 3188
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 5902 3176 5908 3188
rect 5675 3148 5908 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6270 3176 6276 3188
rect 6104 3148 6276 3176
rect 4065 3111 4123 3117
rect 2976 3080 3280 3108
rect 3436 3080 3924 3108
rect 2976 3052 3004 3080
rect 3436 3052 3464 3080
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2866 3040 2872 3052
rect 2547 3012 2872 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 3896 3049 3924 3080
rect 4065 3077 4077 3111
rect 4111 3077 4123 3111
rect 4356 3108 4384 3136
rect 4065 3071 4123 3077
rect 4264 3080 4384 3108
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 2976 2836 3004 3000
rect 3528 2972 3556 3003
rect 3970 3000 3976 3052
rect 4028 3000 4034 3052
rect 4264 3049 4292 3080
rect 4706 3068 4712 3120
rect 4764 3068 4770 3120
rect 4982 3068 4988 3120
rect 5040 3108 5046 3120
rect 5353 3111 5411 3117
rect 5353 3108 5365 3111
rect 5040 3080 5365 3108
rect 5040 3068 5046 3080
rect 5353 3077 5365 3080
rect 5399 3077 5411 3111
rect 5353 3071 5411 3077
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4724 3040 4752 3068
rect 4387 3012 4752 3040
rect 5077 3043 5135 3049
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5166 3040 5172 3052
rect 5123 3012 5172 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5460 3049 5488 3136
rect 5552 3108 5580 3136
rect 5721 3111 5779 3117
rect 5721 3108 5733 3111
rect 5552 3080 5733 3108
rect 5721 3077 5733 3080
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 6104 3049 6132 3148
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7742 3176 7748 3188
rect 7331 3148 7748 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8110 3176 8116 3188
rect 7975 3148 8116 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 8570 3176 8576 3188
rect 8404 3148 8576 3176
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 6656 3108 6684 3136
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 6236 3080 6592 3108
rect 6656 3080 7573 3108
rect 6236 3068 6242 3080
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 3694 2972 3700 2984
rect 3528 2944 3700 2972
rect 3694 2932 3700 2944
rect 3752 2972 3758 2984
rect 3752 2944 4384 2972
rect 3752 2932 3758 2944
rect 4356 2916 4384 2944
rect 4614 2932 4620 2984
rect 4672 2932 4678 2984
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 4948 2944 5212 2972
rect 4948 2932 4954 2944
rect 3786 2904 3792 2916
rect 3436 2876 3792 2904
rect 3436 2845 3464 2876
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 4338 2864 4344 2916
rect 4396 2864 4402 2916
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2904 4583 2907
rect 4632 2904 4660 2932
rect 4571 2876 4660 2904
rect 4571 2873 4583 2876
rect 4525 2867 4583 2873
rect 5074 2864 5080 2916
rect 5132 2864 5138 2916
rect 2823 2808 3004 2836
rect 3421 2839 3479 2845
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3421 2805 3433 2839
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 5092 2836 5120 2864
rect 3743 2808 5120 2836
rect 5184 2836 5212 2944
rect 5276 2904 5304 3003
rect 5920 2972 5948 3003
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 6564 3040 6592 3080
rect 7561 3077 7573 3080
rect 7607 3077 7619 3111
rect 8220 3108 8248 3136
rect 8312 3108 8340 3136
rect 7561 3071 7619 3077
rect 7760 3080 8248 3108
rect 8286 3080 8340 3108
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6564 3012 6745 3040
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 6380 2972 6408 3000
rect 5920 2944 6408 2972
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7392 2972 7420 3003
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7760 3049 7788 3080
rect 8286 3049 8314 3080
rect 8404 3049 8432 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9122 3176 9128 3188
rect 8803 3148 9128 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 12066 3136 12072 3188
rect 12124 3136 12130 3188
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12216 3148 12265 3176
rect 12216 3136 12222 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12526 3136 12532 3188
rect 12584 3136 12590 3188
rect 8481 3111 8539 3117
rect 8481 3077 8493 3111
rect 8527 3108 8539 3111
rect 8662 3108 8668 3120
rect 8527 3080 8668 3108
rect 8527 3077 8539 3080
rect 8481 3071 8539 3077
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8251 3043 8314 3049
rect 8251 3009 8263 3043
rect 8297 3012 8314 3043
rect 8389 3043 8447 3049
rect 8297 3009 8309 3012
rect 8251 3003 8309 3009
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 6687 2944 7512 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6270 2904 6276 2916
rect 5276 2876 6276 2904
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 5184 2808 6469 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 7484 2836 7512 2944
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 8496 2972 8524 3071
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8938 3040 8944 3052
rect 8619 3012 8944 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8076 2944 8524 2972
rect 8076 2932 8082 2944
rect 8588 2836 8616 3003
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9232 3040 9260 3136
rect 9171 3012 9260 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9398 3000 9404 3052
rect 9456 3000 9462 3052
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 12084 3040 12112 3136
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 12084 3012 12173 3040
rect 9493 3003 9551 3009
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 8904 2944 9229 2972
rect 8904 2932 8910 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 7484 2808 8616 2836
rect 9232 2836 9260 2935
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9508 2972 9536 3003
rect 9364 2944 9536 2972
rect 9364 2932 9370 2944
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 12360 2972 12388 3003
rect 12434 3000 12440 3052
rect 12492 3000 12498 3052
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3040 13047 3043
rect 13446 3040 13452 3052
rect 13035 3012 13452 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 10560 2944 12388 2972
rect 10560 2932 10566 2944
rect 9324 2904 9352 2932
rect 9674 2904 9680 2916
rect 9324 2876 9680 2904
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 10928 2876 12817 2904
rect 10928 2864 10934 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 10042 2836 10048 2848
rect 9232 2808 10048 2836
rect 6457 2799 6515 2805
rect 10042 2796 10048 2808
rect 10100 2836 10106 2848
rect 10318 2836 10324 2848
rect 10100 2808 10324 2836
rect 10100 2796 10106 2808
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 1104 2746 13340 2768
rect 1104 2694 2479 2746
rect 2531 2694 2543 2746
rect 2595 2694 2607 2746
rect 2659 2694 2671 2746
rect 2723 2694 2735 2746
rect 2787 2694 5538 2746
rect 5590 2694 5602 2746
rect 5654 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 8597 2746
rect 8649 2694 8661 2746
rect 8713 2694 8725 2746
rect 8777 2694 8789 2746
rect 8841 2694 8853 2746
rect 8905 2694 11656 2746
rect 11708 2694 11720 2746
rect 11772 2694 11784 2746
rect 11836 2694 11848 2746
rect 11900 2694 11912 2746
rect 11964 2694 13340 2746
rect 1104 2672 13340 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 2866 2632 2872 2644
rect 2823 2604 2872 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 2866 2592 2872 2604
rect 2924 2632 2930 2644
rect 3694 2632 3700 2644
rect 2924 2604 3700 2632
rect 2924 2592 2930 2604
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4890 2632 4896 2644
rect 4396 2604 4896 2632
rect 4396 2592 4402 2604
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6086 2632 6092 2644
rect 5951 2604 6092 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6454 2592 6460 2644
rect 6512 2592 6518 2644
rect 8938 2592 8944 2644
rect 8996 2592 9002 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 9732 2604 10425 2632
rect 9732 2592 9738 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 12768 2604 12817 2632
rect 12768 2592 12774 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 6472 2564 6500 2592
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6472 2536 7297 2564
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 6178 2388 6184 2440
rect 6236 2428 6242 2440
rect 6840 2437 6868 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 10376 2468 11805 2496
rect 10376 2456 10382 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6236 2400 6745 2428
rect 6236 2388 6242 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11532 2360 11560 2391
rect 11882 2360 11888 2372
rect 11532 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 12986 2360 12992 2372
rect 12943 2332 12992 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 12986 2320 12992 2332
rect 13044 2320 13050 2372
rect 1104 2202 13499 2224
rect 1104 2150 4008 2202
rect 4060 2150 4072 2202
rect 4124 2150 4136 2202
rect 4188 2150 4200 2202
rect 4252 2150 4264 2202
rect 4316 2150 7067 2202
rect 7119 2150 7131 2202
rect 7183 2150 7195 2202
rect 7247 2150 7259 2202
rect 7311 2150 7323 2202
rect 7375 2150 10126 2202
rect 10178 2150 10190 2202
rect 10242 2150 10254 2202
rect 10306 2150 10318 2202
rect 10370 2150 10382 2202
rect 10434 2150 13185 2202
rect 13237 2150 13249 2202
rect 13301 2150 13313 2202
rect 13365 2150 13377 2202
rect 13429 2150 13441 2202
rect 13493 2150 13499 2202
rect 1104 2128 13499 2150
<< via1 >>
rect 4008 14118 4060 14170
rect 4072 14118 4124 14170
rect 4136 14118 4188 14170
rect 4200 14118 4252 14170
rect 4264 14118 4316 14170
rect 7067 14118 7119 14170
rect 7131 14118 7183 14170
rect 7195 14118 7247 14170
rect 7259 14118 7311 14170
rect 7323 14118 7375 14170
rect 10126 14118 10178 14170
rect 10190 14118 10242 14170
rect 10254 14118 10306 14170
rect 10318 14118 10370 14170
rect 10382 14118 10434 14170
rect 13185 14118 13237 14170
rect 13249 14118 13301 14170
rect 13313 14118 13365 14170
rect 13377 14118 13429 14170
rect 13441 14118 13493 14170
rect 3608 14016 3660 14068
rect 10784 14016 10836 14068
rect 13268 13948 13320 14000
rect 6276 13880 6328 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 12716 13787 12768 13796
rect 12716 13753 12725 13787
rect 12725 13753 12759 13787
rect 12759 13753 12768 13787
rect 12716 13744 12768 13753
rect 2479 13574 2531 13626
rect 2543 13574 2595 13626
rect 2607 13574 2659 13626
rect 2671 13574 2723 13626
rect 2735 13574 2787 13626
rect 5538 13574 5590 13626
rect 5602 13574 5654 13626
rect 5666 13574 5718 13626
rect 5730 13574 5782 13626
rect 5794 13574 5846 13626
rect 8597 13574 8649 13626
rect 8661 13574 8713 13626
rect 8725 13574 8777 13626
rect 8789 13574 8841 13626
rect 8853 13574 8905 13626
rect 11656 13574 11708 13626
rect 11720 13574 11772 13626
rect 11784 13574 11836 13626
rect 11848 13574 11900 13626
rect 11912 13574 11964 13626
rect 6736 13336 6788 13388
rect 6920 13268 6972 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9772 13268 9824 13320
rect 11612 13268 11664 13320
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7748 13132 7800 13184
rect 7840 13132 7892 13184
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 4008 13030 4060 13082
rect 4072 13030 4124 13082
rect 4136 13030 4188 13082
rect 4200 13030 4252 13082
rect 4264 13030 4316 13082
rect 7067 13030 7119 13082
rect 7131 13030 7183 13082
rect 7195 13030 7247 13082
rect 7259 13030 7311 13082
rect 7323 13030 7375 13082
rect 10126 13030 10178 13082
rect 10190 13030 10242 13082
rect 10254 13030 10306 13082
rect 10318 13030 10370 13082
rect 10382 13030 10434 13082
rect 13185 13030 13237 13082
rect 13249 13030 13301 13082
rect 13313 13030 13365 13082
rect 13377 13030 13429 13082
rect 13441 13030 13493 13082
rect 6644 12860 6696 12912
rect 6736 12903 6788 12912
rect 6736 12869 6745 12903
rect 6745 12869 6779 12903
rect 6779 12869 6788 12903
rect 6736 12860 6788 12869
rect 6920 12860 6972 12912
rect 5448 12724 5500 12776
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 6000 12588 6052 12640
rect 7288 12792 7340 12844
rect 9772 12928 9824 12980
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 7840 12860 7892 12912
rect 8484 12860 8536 12912
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 12716 12860 12768 12912
rect 10784 12792 10836 12844
rect 7748 12724 7800 12776
rect 9864 12724 9916 12776
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 10048 12656 10100 12708
rect 8208 12588 8260 12640
rect 10140 12588 10192 12640
rect 2479 12486 2531 12538
rect 2543 12486 2595 12538
rect 2607 12486 2659 12538
rect 2671 12486 2723 12538
rect 2735 12486 2787 12538
rect 5538 12486 5590 12538
rect 5602 12486 5654 12538
rect 5666 12486 5718 12538
rect 5730 12486 5782 12538
rect 5794 12486 5846 12538
rect 8597 12486 8649 12538
rect 8661 12486 8713 12538
rect 8725 12486 8777 12538
rect 8789 12486 8841 12538
rect 8853 12486 8905 12538
rect 11656 12486 11708 12538
rect 11720 12486 11772 12538
rect 11784 12486 11836 12538
rect 11848 12486 11900 12538
rect 11912 12486 11964 12538
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 7288 12384 7340 12436
rect 7472 12384 7524 12436
rect 8116 12384 8168 12436
rect 8484 12384 8536 12436
rect 9128 12384 9180 12436
rect 9772 12384 9824 12436
rect 5080 12248 5132 12257
rect 5632 12112 5684 12164
rect 6000 12112 6052 12164
rect 6736 12112 6788 12164
rect 7380 12248 7432 12300
rect 10784 12384 10836 12436
rect 8208 12248 8260 12300
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9680 12248 9732 12300
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 10048 12316 10100 12368
rect 10140 12316 10192 12368
rect 10232 12316 10284 12368
rect 11980 12384 12032 12436
rect 4068 12044 4120 12096
rect 6368 12044 6420 12096
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 9312 12155 9364 12164
rect 9312 12121 9321 12155
rect 9321 12121 9355 12155
rect 9355 12121 9364 12155
rect 9312 12112 9364 12121
rect 7564 12044 7616 12096
rect 9864 12112 9916 12164
rect 11428 12180 11480 12232
rect 12716 12248 12768 12300
rect 9956 12044 10008 12096
rect 10508 12044 10560 12096
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 4008 11942 4060 11994
rect 4072 11942 4124 11994
rect 4136 11942 4188 11994
rect 4200 11942 4252 11994
rect 4264 11942 4316 11994
rect 7067 11942 7119 11994
rect 7131 11942 7183 11994
rect 7195 11942 7247 11994
rect 7259 11942 7311 11994
rect 7323 11942 7375 11994
rect 10126 11942 10178 11994
rect 10190 11942 10242 11994
rect 10254 11942 10306 11994
rect 10318 11942 10370 11994
rect 10382 11942 10434 11994
rect 13185 11942 13237 11994
rect 13249 11942 13301 11994
rect 13313 11942 13365 11994
rect 13377 11942 13429 11994
rect 13441 11942 13493 11994
rect 6552 11840 6604 11892
rect 9128 11840 9180 11892
rect 10048 11840 10100 11892
rect 11980 11840 12032 11892
rect 5908 11704 5960 11756
rect 7012 11704 7064 11756
rect 6828 11636 6880 11688
rect 6920 11636 6972 11688
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 9496 11636 9548 11688
rect 10140 11747 10192 11756
rect 10140 11713 10150 11747
rect 10150 11713 10184 11747
rect 10184 11713 10192 11747
rect 10140 11704 10192 11713
rect 10324 11704 10376 11756
rect 10508 11704 10560 11756
rect 11152 11679 11204 11688
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 11520 11636 11572 11688
rect 9772 11611 9824 11620
rect 9772 11577 9781 11611
rect 9781 11577 9815 11611
rect 9815 11577 9824 11611
rect 9772 11568 9824 11577
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 7196 11500 7248 11552
rect 8024 11500 8076 11552
rect 9404 11500 9456 11552
rect 10232 11500 10284 11552
rect 10692 11500 10744 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11336 11500 11388 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 2479 11398 2531 11450
rect 2543 11398 2595 11450
rect 2607 11398 2659 11450
rect 2671 11398 2723 11450
rect 2735 11398 2787 11450
rect 5538 11398 5590 11450
rect 5602 11398 5654 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 8597 11398 8649 11450
rect 8661 11398 8713 11450
rect 8725 11398 8777 11450
rect 8789 11398 8841 11450
rect 8853 11398 8905 11450
rect 11656 11398 11708 11450
rect 11720 11398 11772 11450
rect 11784 11398 11836 11450
rect 11848 11398 11900 11450
rect 11912 11398 11964 11450
rect 4620 11296 4672 11348
rect 6644 11296 6696 11348
rect 6920 11296 6972 11348
rect 7012 11228 7064 11280
rect 7564 11296 7616 11348
rect 9312 11296 9364 11348
rect 9956 11296 10008 11348
rect 11060 11296 11112 11348
rect 11152 11339 11204 11348
rect 11152 11305 11161 11339
rect 11161 11305 11195 11339
rect 11195 11305 11204 11339
rect 11152 11296 11204 11305
rect 11428 11296 11480 11348
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 5080 11092 5132 11144
rect 4712 11024 4764 11076
rect 6920 11092 6972 11144
rect 7748 11092 7800 11144
rect 9772 11160 9824 11212
rect 10876 11160 10928 11212
rect 8024 11024 8076 11076
rect 8392 11024 8444 11076
rect 6644 10956 6696 11008
rect 7196 10956 7248 11008
rect 9404 11092 9456 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 10508 11092 10560 11144
rect 11152 11024 11204 11076
rect 11336 11092 11388 11144
rect 11520 11092 11572 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 12256 11092 12308 11144
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 10048 10956 10100 11008
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 4008 10854 4060 10906
rect 4072 10854 4124 10906
rect 4136 10854 4188 10906
rect 4200 10854 4252 10906
rect 4264 10854 4316 10906
rect 7067 10854 7119 10906
rect 7131 10854 7183 10906
rect 7195 10854 7247 10906
rect 7259 10854 7311 10906
rect 7323 10854 7375 10906
rect 10126 10854 10178 10906
rect 10190 10854 10242 10906
rect 10254 10854 10306 10906
rect 10318 10854 10370 10906
rect 10382 10854 10434 10906
rect 13185 10854 13237 10906
rect 13249 10854 13301 10906
rect 13313 10854 13365 10906
rect 13377 10854 13429 10906
rect 13441 10854 13493 10906
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 5448 10752 5500 10804
rect 5908 10752 5960 10804
rect 6644 10684 6696 10736
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 7012 10616 7064 10668
rect 7748 10616 7800 10668
rect 8024 10616 8076 10668
rect 6736 10480 6788 10532
rect 7104 10548 7156 10600
rect 9496 10752 9548 10804
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 11152 10752 11204 10804
rect 8392 10727 8444 10736
rect 8392 10693 8401 10727
rect 8401 10693 8435 10727
rect 8435 10693 8444 10727
rect 8392 10684 8444 10693
rect 9680 10684 9732 10736
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10140 10548 10192 10600
rect 10600 10480 10652 10532
rect 11520 10616 11572 10668
rect 11980 10752 12032 10804
rect 11060 10548 11112 10600
rect 12624 10548 12676 10600
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 11520 10523 11572 10532
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 11520 10489 11529 10523
rect 11529 10489 11563 10523
rect 11563 10489 11572 10523
rect 11520 10480 11572 10489
rect 11796 10480 11848 10532
rect 12256 10480 12308 10532
rect 11428 10412 11480 10464
rect 11980 10412 12032 10464
rect 2479 10310 2531 10362
rect 2543 10310 2595 10362
rect 2607 10310 2659 10362
rect 2671 10310 2723 10362
rect 2735 10310 2787 10362
rect 5538 10310 5590 10362
rect 5602 10310 5654 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 8597 10310 8649 10362
rect 8661 10310 8713 10362
rect 8725 10310 8777 10362
rect 8789 10310 8841 10362
rect 8853 10310 8905 10362
rect 11656 10310 11708 10362
rect 11720 10310 11772 10362
rect 11784 10310 11836 10362
rect 11848 10310 11900 10362
rect 11912 10310 11964 10362
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 9404 10208 9456 10260
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 10600 10208 10652 10260
rect 11520 10208 11572 10260
rect 11980 10208 12032 10260
rect 12164 10208 12216 10260
rect 12716 10208 12768 10260
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5908 10072 5960 10124
rect 7104 10072 7156 10124
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 6000 9936 6052 9988
rect 10048 9936 10100 9988
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 7748 9868 7800 9920
rect 9956 9868 10008 9920
rect 11244 10004 11296 10056
rect 11520 10047 11572 10056
rect 11520 10013 11530 10047
rect 11530 10013 11564 10047
rect 11564 10013 11572 10047
rect 11520 10004 11572 10013
rect 12072 10004 12124 10056
rect 12256 10004 12308 10056
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 4008 9766 4060 9818
rect 4072 9766 4124 9818
rect 4136 9766 4188 9818
rect 4200 9766 4252 9818
rect 4264 9766 4316 9818
rect 7067 9766 7119 9818
rect 7131 9766 7183 9818
rect 7195 9766 7247 9818
rect 7259 9766 7311 9818
rect 7323 9766 7375 9818
rect 10126 9766 10178 9818
rect 10190 9766 10242 9818
rect 10254 9766 10306 9818
rect 10318 9766 10370 9818
rect 10382 9766 10434 9818
rect 13185 9766 13237 9818
rect 13249 9766 13301 9818
rect 13313 9766 13365 9818
rect 13377 9766 13429 9818
rect 13441 9766 13493 9818
rect 5448 9664 5500 9716
rect 3148 9596 3200 9648
rect 6000 9707 6052 9716
rect 6000 9673 6009 9707
rect 6009 9673 6043 9707
rect 6043 9673 6052 9707
rect 6000 9664 6052 9673
rect 7472 9664 7524 9716
rect 8208 9664 8260 9716
rect 11520 9664 11572 9716
rect 11612 9707 11664 9716
rect 11612 9673 11621 9707
rect 11621 9673 11655 9707
rect 11655 9673 11664 9707
rect 11612 9664 11664 9673
rect 3240 9324 3292 9376
rect 3424 9324 3476 9376
rect 7564 9528 7616 9580
rect 8484 9596 8536 9648
rect 10508 9596 10560 9648
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 10048 9528 10100 9580
rect 10692 9528 10744 9580
rect 11152 9596 11204 9648
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 10968 9528 11020 9580
rect 11428 9528 11480 9580
rect 12716 9528 12768 9580
rect 10876 9392 10928 9444
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 10692 9324 10744 9376
rect 12624 9324 12676 9376
rect 2479 9222 2531 9274
rect 2543 9222 2595 9274
rect 2607 9222 2659 9274
rect 2671 9222 2723 9274
rect 2735 9222 2787 9274
rect 5538 9222 5590 9274
rect 5602 9222 5654 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 8597 9222 8649 9274
rect 8661 9222 8713 9274
rect 8725 9222 8777 9274
rect 8789 9222 8841 9274
rect 8853 9222 8905 9274
rect 11656 9222 11708 9274
rect 11720 9222 11772 9274
rect 11784 9222 11836 9274
rect 11848 9222 11900 9274
rect 11912 9222 11964 9274
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 5080 8984 5132 9036
rect 5172 8984 5224 9036
rect 7748 9120 7800 9172
rect 3424 8916 3476 8968
rect 4344 8916 4396 8968
rect 6092 8984 6144 9036
rect 8484 9120 8536 9172
rect 11520 9052 11572 9104
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 7380 8916 7432 8968
rect 7564 8916 7616 8968
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2964 8891 3016 8900
rect 2964 8857 2973 8891
rect 2973 8857 3007 8891
rect 3007 8857 3016 8891
rect 2964 8848 3016 8857
rect 3792 8848 3844 8900
rect 3884 8780 3936 8832
rect 5172 8848 5224 8900
rect 5724 8891 5776 8900
rect 5724 8857 5733 8891
rect 5733 8857 5767 8891
rect 5767 8857 5776 8891
rect 5724 8848 5776 8857
rect 12348 9120 12400 9172
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 4528 8780 4580 8832
rect 8300 8780 8352 8832
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 4008 8678 4060 8730
rect 4072 8678 4124 8730
rect 4136 8678 4188 8730
rect 4200 8678 4252 8730
rect 4264 8678 4316 8730
rect 7067 8678 7119 8730
rect 7131 8678 7183 8730
rect 7195 8678 7247 8730
rect 7259 8678 7311 8730
rect 7323 8678 7375 8730
rect 10126 8678 10178 8730
rect 10190 8678 10242 8730
rect 10254 8678 10306 8730
rect 10318 8678 10370 8730
rect 10382 8678 10434 8730
rect 13185 8678 13237 8730
rect 13249 8678 13301 8730
rect 13313 8678 13365 8730
rect 13377 8678 13429 8730
rect 13441 8678 13493 8730
rect 1492 8576 1544 8628
rect 2044 8576 2096 8628
rect 2964 8576 3016 8628
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 3332 8576 3384 8585
rect 4344 8576 4396 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 12348 8619 12400 8628
rect 12348 8585 12357 8619
rect 12357 8585 12391 8619
rect 12391 8585 12400 8619
rect 12348 8576 12400 8585
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3332 8440 3384 8492
rect 3792 8440 3844 8492
rect 4620 8508 4672 8560
rect 5172 8508 5224 8560
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 6368 8551 6420 8560
rect 6368 8517 6377 8551
rect 6377 8517 6411 8551
rect 6411 8517 6420 8551
rect 6368 8508 6420 8517
rect 2412 8372 2464 8424
rect 8024 8440 8076 8492
rect 8208 8440 8260 8492
rect 10508 8440 10560 8492
rect 12256 8440 12308 8492
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 3884 8347 3936 8356
rect 3884 8313 3893 8347
rect 3893 8313 3927 8347
rect 3927 8313 3936 8347
rect 3884 8304 3936 8313
rect 2780 8236 2832 8288
rect 2964 8236 3016 8288
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 2479 8134 2531 8186
rect 2543 8134 2595 8186
rect 2607 8134 2659 8186
rect 2671 8134 2723 8186
rect 2735 8134 2787 8186
rect 5538 8134 5590 8186
rect 5602 8134 5654 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 8597 8134 8649 8186
rect 8661 8134 8713 8186
rect 8725 8134 8777 8186
rect 8789 8134 8841 8186
rect 8853 8134 8905 8186
rect 11656 8134 11708 8186
rect 11720 8134 11772 8186
rect 11784 8134 11836 8186
rect 11848 8134 11900 8186
rect 11912 8134 11964 8186
rect 2872 8032 2924 8084
rect 3792 8032 3844 8084
rect 5080 8032 5132 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 2780 7964 2832 8016
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 2320 7760 2372 7812
rect 3148 7828 3200 7880
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 4344 7828 4396 7880
rect 6644 7828 6696 7880
rect 7656 7828 7708 7880
rect 8484 7828 8536 7880
rect 9220 7828 9272 7880
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 8944 7803 8996 7812
rect 8944 7769 8953 7803
rect 8953 7769 8987 7803
rect 8987 7769 8996 7803
rect 8944 7760 8996 7769
rect 9404 7760 9456 7812
rect 12164 7760 12216 7812
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 8300 7692 8352 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 4008 7590 4060 7642
rect 4072 7590 4124 7642
rect 4136 7590 4188 7642
rect 4200 7590 4252 7642
rect 4264 7590 4316 7642
rect 7067 7590 7119 7642
rect 7131 7590 7183 7642
rect 7195 7590 7247 7642
rect 7259 7590 7311 7642
rect 7323 7590 7375 7642
rect 10126 7590 10178 7642
rect 10190 7590 10242 7642
rect 10254 7590 10306 7642
rect 10318 7590 10370 7642
rect 10382 7590 10434 7642
rect 13185 7590 13237 7642
rect 13249 7590 13301 7642
rect 13313 7590 13365 7642
rect 13377 7590 13429 7642
rect 13441 7590 13493 7642
rect 2412 7488 2464 7540
rect 8392 7488 8444 7540
rect 6092 7420 6144 7472
rect 8024 7420 8076 7472
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 2320 7352 2372 7404
rect 3148 7352 3200 7404
rect 4988 7216 5040 7268
rect 9036 7395 9088 7404
rect 9036 7361 9056 7395
rect 9056 7361 9088 7395
rect 9036 7352 9088 7361
rect 12256 7284 12308 7336
rect 6184 7216 6236 7268
rect 2780 7148 2832 7200
rect 4804 7148 4856 7200
rect 5816 7148 5868 7200
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 6552 7148 6604 7200
rect 7564 7148 7616 7200
rect 9496 7148 9548 7200
rect 10140 7148 10192 7200
rect 12164 7148 12216 7200
rect 2479 7046 2531 7098
rect 2543 7046 2595 7098
rect 2607 7046 2659 7098
rect 2671 7046 2723 7098
rect 2735 7046 2787 7098
rect 5538 7046 5590 7098
rect 5602 7046 5654 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 8597 7046 8649 7098
rect 8661 7046 8713 7098
rect 8725 7046 8777 7098
rect 8789 7046 8841 7098
rect 8853 7046 8905 7098
rect 11656 7046 11708 7098
rect 11720 7046 11772 7098
rect 11784 7046 11836 7098
rect 11848 7046 11900 7098
rect 11912 7046 11964 7098
rect 2228 6944 2280 6996
rect 5908 6944 5960 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 5448 6808 5500 6860
rect 5908 6808 5960 6860
rect 8484 6944 8536 6996
rect 9220 6944 9272 6996
rect 9588 6944 9640 6996
rect 10784 6944 10836 6996
rect 11152 6851 11204 6860
rect 2964 6740 3016 6792
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 3700 6672 3752 6724
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 4436 6672 4488 6724
rect 5356 6672 5408 6724
rect 6092 6672 6144 6724
rect 6552 6672 6604 6724
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 4712 6647 4764 6656
rect 4712 6613 4721 6647
rect 4721 6613 4755 6647
rect 4755 6613 4764 6647
rect 4712 6604 4764 6613
rect 8944 6740 8996 6792
rect 9036 6740 9088 6792
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 9772 6740 9824 6792
rect 9864 6740 9916 6792
rect 9312 6715 9364 6724
rect 9312 6681 9321 6715
rect 9321 6681 9355 6715
rect 9355 6681 9364 6715
rect 9312 6672 9364 6681
rect 7656 6604 7708 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 10048 6604 10100 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 12164 6672 12216 6724
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 4008 6502 4060 6554
rect 4072 6502 4124 6554
rect 4136 6502 4188 6554
rect 4200 6502 4252 6554
rect 4264 6502 4316 6554
rect 7067 6502 7119 6554
rect 7131 6502 7183 6554
rect 7195 6502 7247 6554
rect 7259 6502 7311 6554
rect 7323 6502 7375 6554
rect 10126 6502 10178 6554
rect 10190 6502 10242 6554
rect 10254 6502 10306 6554
rect 10318 6502 10370 6554
rect 10382 6502 10434 6554
rect 13185 6502 13237 6554
rect 13249 6502 13301 6554
rect 13313 6502 13365 6554
rect 13377 6502 13429 6554
rect 13441 6502 13493 6554
rect 4436 6400 4488 6452
rect 4712 6400 4764 6452
rect 4988 6400 5040 6452
rect 7656 6400 7708 6452
rect 2964 6264 3016 6316
rect 3884 6264 3936 6316
rect 3056 6196 3108 6248
rect 4344 6332 4396 6384
rect 5908 6332 5960 6384
rect 7564 6332 7616 6384
rect 8392 6400 8444 6452
rect 9496 6443 9548 6452
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 9772 6400 9824 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10600 6400 10652 6452
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 10048 6264 10100 6316
rect 4344 6239 4396 6248
rect 4344 6205 4360 6239
rect 4360 6205 4394 6239
rect 4394 6205 4396 6239
rect 4344 6196 4396 6205
rect 5264 6196 5316 6248
rect 9772 6196 9824 6248
rect 12900 6332 12952 6384
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 2136 6060 2188 6112
rect 2872 6060 2924 6112
rect 3332 6060 3384 6112
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 3792 6060 3844 6112
rect 4344 6060 4396 6112
rect 4804 6060 4856 6112
rect 6184 6060 6236 6112
rect 8300 6060 8352 6112
rect 2479 5958 2531 6010
rect 2543 5958 2595 6010
rect 2607 5958 2659 6010
rect 2671 5958 2723 6010
rect 2735 5958 2787 6010
rect 5538 5958 5590 6010
rect 5602 5958 5654 6010
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 8597 5958 8649 6010
rect 8661 5958 8713 6010
rect 8725 5958 8777 6010
rect 8789 5958 8841 6010
rect 8853 5958 8905 6010
rect 11656 5958 11708 6010
rect 11720 5958 11772 6010
rect 11784 5958 11836 6010
rect 11848 5958 11900 6010
rect 11912 5958 11964 6010
rect 1400 5720 1452 5772
rect 4252 5856 4304 5908
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 4896 5856 4948 5908
rect 6276 5856 6328 5908
rect 7472 5856 7524 5908
rect 8760 5856 8812 5908
rect 2136 5720 2188 5772
rect 4436 5720 4488 5772
rect 4528 5720 4580 5772
rect 5448 5788 5500 5840
rect 9036 5720 9088 5772
rect 2872 5652 2924 5704
rect 6644 5652 6696 5704
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 3700 5516 3752 5568
rect 4008 5414 4060 5466
rect 4072 5414 4124 5466
rect 4136 5414 4188 5466
rect 4200 5414 4252 5466
rect 4264 5414 4316 5466
rect 7067 5414 7119 5466
rect 7131 5414 7183 5466
rect 7195 5414 7247 5466
rect 7259 5414 7311 5466
rect 7323 5414 7375 5466
rect 10126 5414 10178 5466
rect 10190 5414 10242 5466
rect 10254 5414 10306 5466
rect 10318 5414 10370 5466
rect 10382 5414 10434 5466
rect 13185 5414 13237 5466
rect 13249 5414 13301 5466
rect 13313 5414 13365 5466
rect 13377 5414 13429 5466
rect 13441 5414 13493 5466
rect 3056 5312 3108 5364
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 5264 5312 5316 5364
rect 5908 5312 5960 5364
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 9496 5312 9548 5364
rect 9772 5312 9824 5364
rect 9864 5312 9916 5364
rect 3884 5244 3936 5296
rect 5540 5287 5592 5296
rect 5540 5253 5549 5287
rect 5549 5253 5583 5287
rect 5583 5253 5592 5287
rect 5540 5244 5592 5253
rect 6920 5244 6972 5296
rect 8300 5287 8352 5296
rect 8300 5253 8317 5287
rect 8317 5253 8352 5287
rect 8300 5244 8352 5253
rect 9128 5244 9180 5296
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 3700 5176 3752 5228
rect 2964 5108 3016 5160
rect 6092 5176 6144 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9220 5176 9272 5228
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10784 5176 10836 5228
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 11244 5108 11296 5160
rect 5172 5040 5224 5092
rect 12440 5108 12492 5160
rect 2136 4972 2188 5024
rect 4344 4972 4396 5024
rect 9404 4972 9456 5024
rect 9772 4972 9824 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 12164 4972 12216 5024
rect 2479 4870 2531 4922
rect 2543 4870 2595 4922
rect 2607 4870 2659 4922
rect 2671 4870 2723 4922
rect 2735 4870 2787 4922
rect 5538 4870 5590 4922
rect 5602 4870 5654 4922
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 8597 4870 8649 4922
rect 8661 4870 8713 4922
rect 8725 4870 8777 4922
rect 8789 4870 8841 4922
rect 8853 4870 8905 4922
rect 11656 4870 11708 4922
rect 11720 4870 11772 4922
rect 11784 4870 11836 4922
rect 11848 4870 11900 4922
rect 11912 4870 11964 4922
rect 9220 4768 9272 4820
rect 5172 4632 5224 4684
rect 11520 4632 11572 4684
rect 940 4564 992 4616
rect 2136 4564 2188 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 10968 4496 11020 4548
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 12164 4496 12216 4548
rect 11060 4428 11112 4480
rect 11336 4428 11388 4480
rect 4008 4326 4060 4378
rect 4072 4326 4124 4378
rect 4136 4326 4188 4378
rect 4200 4326 4252 4378
rect 4264 4326 4316 4378
rect 7067 4326 7119 4378
rect 7131 4326 7183 4378
rect 7195 4326 7247 4378
rect 7259 4326 7311 4378
rect 7323 4326 7375 4378
rect 10126 4326 10178 4378
rect 10190 4326 10242 4378
rect 10254 4326 10306 4378
rect 10318 4326 10370 4378
rect 10382 4326 10434 4378
rect 13185 4326 13237 4378
rect 13249 4326 13301 4378
rect 13313 4326 13365 4378
rect 13377 4326 13429 4378
rect 13441 4326 13493 4378
rect 3608 4224 3660 4276
rect 2320 4088 2372 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 4068 4156 4120 4208
rect 2044 4020 2096 4072
rect 3148 3952 3200 4004
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 4988 4088 5040 4140
rect 6092 4088 6144 4140
rect 7656 4224 7708 4276
rect 8484 4224 8536 4276
rect 10784 4224 10836 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 11336 4224 11388 4276
rect 7288 4088 7340 4140
rect 2872 3884 2924 3936
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 3056 3884 3108 3936
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 4068 3995 4120 4004
rect 4068 3961 4077 3995
rect 4077 3961 4111 3995
rect 4111 3961 4120 3995
rect 4068 3952 4120 3961
rect 4252 3952 4304 4004
rect 4712 3952 4764 4004
rect 3700 3884 3752 3936
rect 3792 3884 3844 3936
rect 4344 3884 4396 3936
rect 5080 3884 5132 3936
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 5908 4020 5960 4072
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6644 4020 6696 4072
rect 6828 4020 6880 4072
rect 7104 3995 7156 4004
rect 7104 3961 7113 3995
rect 7113 3961 7147 3995
rect 7147 3961 7156 3995
rect 7104 3952 7156 3961
rect 6644 3884 6696 3936
rect 6736 3884 6788 3936
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 8116 4088 8168 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 7656 3952 7708 4004
rect 9128 4156 9180 4208
rect 9036 4088 9088 4140
rect 9772 4088 9824 4140
rect 11060 4156 11112 4208
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 8760 3884 8812 3936
rect 8944 3884 8996 3936
rect 9036 3884 9088 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 10508 3952 10560 4004
rect 11244 4020 11296 4072
rect 10784 3884 10836 3936
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 2479 3782 2531 3834
rect 2543 3782 2595 3834
rect 2607 3782 2659 3834
rect 2671 3782 2723 3834
rect 2735 3782 2787 3834
rect 5538 3782 5590 3834
rect 5602 3782 5654 3834
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 8597 3782 8649 3834
rect 8661 3782 8713 3834
rect 8725 3782 8777 3834
rect 8789 3782 8841 3834
rect 8853 3782 8905 3834
rect 11656 3782 11708 3834
rect 11720 3782 11772 3834
rect 11784 3782 11836 3834
rect 11848 3782 11900 3834
rect 11912 3782 11964 3834
rect 1584 3544 1636 3596
rect 2228 3612 2280 3664
rect 2044 3544 2096 3596
rect 2872 3680 2924 3732
rect 3148 3544 3200 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3332 3612 3384 3664
rect 3884 3612 3936 3664
rect 4804 3680 4856 3732
rect 5080 3680 5132 3732
rect 6828 3680 6880 3732
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 7104 3680 7156 3732
rect 8024 3680 8076 3732
rect 3608 3476 3660 3528
rect 5448 3612 5500 3664
rect 4252 3476 4304 3528
rect 2044 3340 2096 3392
rect 2872 3383 2924 3392
rect 2872 3349 2881 3383
rect 2881 3349 2915 3383
rect 2915 3349 2924 3383
rect 2872 3340 2924 3349
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 5264 3476 5316 3528
rect 6092 3612 6144 3664
rect 7748 3612 7800 3664
rect 7840 3612 7892 3664
rect 9312 3680 9364 3732
rect 10048 3680 10100 3732
rect 10692 3680 10744 3732
rect 10876 3680 10928 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 6000 3544 6052 3596
rect 6276 3544 6328 3596
rect 6736 3544 6788 3596
rect 6920 3544 6972 3596
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 6368 3476 6420 3528
rect 7288 3476 7340 3528
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8668 3544 8720 3596
rect 8944 3544 8996 3596
rect 9036 3544 9088 3596
rect 6920 3451 6972 3460
rect 6920 3417 6929 3451
rect 6929 3417 6963 3451
rect 6963 3417 6972 3451
rect 6920 3408 6972 3417
rect 5540 3340 5592 3392
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 7748 3340 7800 3392
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 8300 3340 8352 3392
rect 8576 3451 8628 3460
rect 8576 3417 8585 3451
rect 8585 3417 8619 3451
rect 8619 3417 8628 3451
rect 8576 3408 8628 3417
rect 8852 3408 8904 3460
rect 9772 3612 9824 3664
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9404 3476 9456 3528
rect 9680 3519 9732 3528
rect 9680 3485 9690 3519
rect 9690 3485 9724 3519
rect 9724 3485 9732 3519
rect 9680 3476 9732 3485
rect 9772 3476 9824 3528
rect 10048 3519 10100 3528
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 10048 3485 10062 3519
rect 10062 3485 10096 3519
rect 10096 3485 10100 3519
rect 10048 3476 10100 3485
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 10968 3476 11020 3528
rect 12532 3476 12584 3528
rect 9404 3340 9456 3392
rect 12164 3340 12216 3392
rect 4008 3238 4060 3290
rect 4072 3238 4124 3290
rect 4136 3238 4188 3290
rect 4200 3238 4252 3290
rect 4264 3238 4316 3290
rect 7067 3238 7119 3290
rect 7131 3238 7183 3290
rect 7195 3238 7247 3290
rect 7259 3238 7311 3290
rect 7323 3238 7375 3290
rect 10126 3238 10178 3290
rect 10190 3238 10242 3290
rect 10254 3238 10306 3290
rect 10318 3238 10370 3290
rect 10382 3238 10434 3290
rect 13185 3238 13237 3290
rect 13249 3238 13301 3290
rect 13313 3238 13365 3290
rect 13377 3238 13429 3290
rect 13441 3238 13493 3290
rect 2872 3136 2924 3188
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 4252 3136 4304 3188
rect 4344 3136 4396 3188
rect 4896 3136 4948 3188
rect 5448 3136 5500 3188
rect 5540 3136 5592 3188
rect 5908 3136 5960 3188
rect 2872 3000 2924 3052
rect 2964 3000 3016 3052
rect 3424 3000 3476 3052
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4712 3068 4764 3120
rect 4988 3068 5040 3120
rect 5172 3000 5224 3052
rect 6276 3136 6328 3188
rect 6644 3136 6696 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 7748 3136 7800 3188
rect 8116 3136 8168 3188
rect 8208 3136 8260 3188
rect 8300 3136 8352 3188
rect 6184 3068 6236 3120
rect 3700 2932 3752 2984
rect 4620 2932 4672 2984
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 3792 2864 3844 2916
rect 4344 2864 4396 2916
rect 5080 2864 5132 2916
rect 6368 3000 6420 3052
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8576 3136 8628 3188
rect 9128 3136 9180 3188
rect 9220 3136 9272 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 12072 3136 12124 3188
rect 12164 3136 12216 3188
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 6276 2864 6328 2916
rect 8024 2932 8076 2984
rect 8668 3068 8720 3120
rect 8944 3000 8996 3052
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 8852 2932 8904 2984
rect 9312 2932 9364 2984
rect 10508 2932 10560 2984
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 13452 3000 13504 3052
rect 9680 2864 9732 2916
rect 10876 2864 10928 2916
rect 10048 2796 10100 2848
rect 10324 2796 10376 2848
rect 2479 2694 2531 2746
rect 2543 2694 2595 2746
rect 2607 2694 2659 2746
rect 2671 2694 2723 2746
rect 2735 2694 2787 2746
rect 5538 2694 5590 2746
rect 5602 2694 5654 2746
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 8597 2694 8649 2746
rect 8661 2694 8713 2746
rect 8725 2694 8777 2746
rect 8789 2694 8841 2746
rect 8853 2694 8905 2746
rect 11656 2694 11708 2746
rect 11720 2694 11772 2746
rect 11784 2694 11836 2746
rect 11848 2694 11900 2746
rect 11912 2694 11964 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2872 2592 2924 2644
rect 3700 2592 3752 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4896 2592 4948 2644
rect 6092 2592 6144 2644
rect 6460 2592 6512 2644
rect 8944 2635 8996 2644
rect 8944 2601 8953 2635
rect 8953 2601 8987 2635
rect 8987 2601 8996 2635
rect 8944 2592 8996 2601
rect 9680 2592 9732 2644
rect 12716 2592 12768 2644
rect 940 2388 992 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6184 2388 6236 2440
rect 10324 2456 10376 2508
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8760 2388 8812 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11888 2320 11940 2372
rect 12992 2320 13044 2372
rect 4008 2150 4060 2202
rect 4072 2150 4124 2202
rect 4136 2150 4188 2202
rect 4200 2150 4252 2202
rect 4264 2150 4316 2202
rect 7067 2150 7119 2202
rect 7131 2150 7183 2202
rect 7195 2150 7247 2202
rect 7259 2150 7311 2202
rect 7323 2150 7375 2202
rect 10126 2150 10178 2202
rect 10190 2150 10242 2202
rect 10254 2150 10306 2202
rect 10318 2150 10370 2202
rect 10382 2150 10434 2202
rect 13185 2150 13237 2202
rect 13249 2150 13301 2202
rect 13313 2150 13365 2202
rect 13377 2150 13429 2202
rect 13441 2150 13493 2202
<< metal2 >>
rect 3606 15801 3662 16601
rect 10782 15801 10838 16601
rect 3620 14074 3648 15801
rect 4008 14172 4316 14181
rect 4008 14170 4014 14172
rect 4070 14170 4094 14172
rect 4150 14170 4174 14172
rect 4230 14170 4254 14172
rect 4310 14170 4316 14172
rect 4070 14118 4072 14170
rect 4252 14118 4254 14170
rect 4008 14116 4014 14118
rect 4070 14116 4094 14118
rect 4150 14116 4174 14118
rect 4230 14116 4254 14118
rect 4310 14116 4316 14118
rect 4008 14107 4316 14116
rect 7067 14172 7375 14181
rect 7067 14170 7073 14172
rect 7129 14170 7153 14172
rect 7209 14170 7233 14172
rect 7289 14170 7313 14172
rect 7369 14170 7375 14172
rect 7129 14118 7131 14170
rect 7311 14118 7313 14170
rect 7067 14116 7073 14118
rect 7129 14116 7153 14118
rect 7209 14116 7233 14118
rect 7289 14116 7313 14118
rect 7369 14116 7375 14118
rect 7067 14107 7375 14116
rect 10126 14172 10434 14181
rect 10126 14170 10132 14172
rect 10188 14170 10212 14172
rect 10268 14170 10292 14172
rect 10348 14170 10372 14172
rect 10428 14170 10434 14172
rect 10188 14118 10190 14170
rect 10370 14118 10372 14170
rect 10126 14116 10132 14118
rect 10188 14116 10212 14118
rect 10268 14116 10292 14118
rect 10348 14116 10372 14118
rect 10428 14116 10434 14118
rect 10126 14107 10434 14116
rect 10796 14074 10824 15801
rect 13185 14172 13493 14181
rect 13185 14170 13191 14172
rect 13247 14170 13271 14172
rect 13327 14170 13351 14172
rect 13407 14170 13431 14172
rect 13487 14170 13493 14172
rect 13247 14118 13249 14170
rect 13429 14118 13431 14170
rect 13185 14116 13191 14118
rect 13247 14116 13271 14118
rect 13327 14116 13351 14118
rect 13407 14116 13431 14118
rect 13487 14116 13493 14118
rect 13185 14107 13493 14116
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 13268 14000 13320 14006
rect 13266 13968 13268 13977
rect 13320 13968 13322 13977
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 10968 13932 11020 13938
rect 13266 13903 13322 13912
rect 10968 13874 11020 13880
rect 2479 13628 2787 13637
rect 2479 13626 2485 13628
rect 2541 13626 2565 13628
rect 2621 13626 2645 13628
rect 2701 13626 2725 13628
rect 2781 13626 2787 13628
rect 2541 13574 2543 13626
rect 2723 13574 2725 13626
rect 2479 13572 2485 13574
rect 2541 13572 2565 13574
rect 2621 13572 2645 13574
rect 2701 13572 2725 13574
rect 2781 13572 2787 13574
rect 2479 13563 2787 13572
rect 5538 13628 5846 13637
rect 5538 13626 5544 13628
rect 5600 13626 5624 13628
rect 5680 13626 5704 13628
rect 5760 13626 5784 13628
rect 5840 13626 5846 13628
rect 5600 13574 5602 13626
rect 5782 13574 5784 13626
rect 5538 13572 5544 13574
rect 5600 13572 5624 13574
rect 5680 13572 5704 13574
rect 5760 13572 5784 13574
rect 5840 13572 5846 13574
rect 5538 13563 5846 13572
rect 4008 13084 4316 13093
rect 4008 13082 4014 13084
rect 4070 13082 4094 13084
rect 4150 13082 4174 13084
rect 4230 13082 4254 13084
rect 4310 13082 4316 13084
rect 4070 13030 4072 13082
rect 4252 13030 4254 13082
rect 4008 13028 4014 13030
rect 4070 13028 4094 13030
rect 4150 13028 4174 13030
rect 4230 13028 4254 13030
rect 4310 13028 4316 13030
rect 4008 13019 4316 13028
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 2479 12540 2787 12549
rect 2479 12538 2485 12540
rect 2541 12538 2565 12540
rect 2621 12538 2645 12540
rect 2701 12538 2725 12540
rect 2781 12538 2787 12540
rect 2541 12486 2543 12538
rect 2723 12486 2725 12538
rect 2479 12484 2485 12486
rect 2541 12484 2565 12486
rect 2621 12484 2645 12486
rect 2701 12484 2725 12486
rect 2781 12484 2787 12486
rect 2479 12475 2787 12484
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 5080 12300 5132 12306
rect 4080 12102 4108 12271
rect 5080 12242 5132 12248
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4008 11996 4316 12005
rect 4008 11994 4014 11996
rect 4070 11994 4094 11996
rect 4150 11994 4174 11996
rect 4230 11994 4254 11996
rect 4310 11994 4316 11996
rect 4070 11942 4072 11994
rect 4252 11942 4254 11994
rect 4008 11940 4014 11942
rect 4070 11940 4094 11942
rect 4150 11940 4174 11942
rect 4230 11940 4254 11942
rect 4310 11940 4316 11942
rect 4008 11931 4316 11940
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 2479 11452 2787 11461
rect 2479 11450 2485 11452
rect 2541 11450 2565 11452
rect 2621 11450 2645 11452
rect 2701 11450 2725 11452
rect 2781 11450 2787 11452
rect 2541 11398 2543 11450
rect 2723 11398 2725 11450
rect 2479 11396 2485 11398
rect 2541 11396 2565 11398
rect 2621 11396 2645 11398
rect 2701 11396 2725 11398
rect 2781 11396 2787 11398
rect 2479 11387 2787 11396
rect 4632 11354 4660 11494
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 5092 11150 5120 12242
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4008 10908 4316 10917
rect 4008 10906 4014 10908
rect 4070 10906 4094 10908
rect 4150 10906 4174 10908
rect 4230 10906 4254 10908
rect 4310 10906 4316 10908
rect 4070 10854 4072 10906
rect 4252 10854 4254 10906
rect 4008 10852 4014 10854
rect 4070 10852 4094 10854
rect 4150 10852 4174 10854
rect 4230 10852 4254 10854
rect 4310 10852 4316 10854
rect 4008 10843 4316 10852
rect 4724 10810 4752 11018
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 2479 10364 2787 10373
rect 2479 10362 2485 10364
rect 2541 10362 2565 10364
rect 2621 10362 2645 10364
rect 2701 10362 2725 10364
rect 2781 10362 2787 10364
rect 2541 10310 2543 10362
rect 2723 10310 2725 10362
rect 2479 10308 2485 10310
rect 2541 10308 2565 10310
rect 2621 10308 2645 10310
rect 2701 10308 2725 10310
rect 2781 10308 2787 10310
rect 2479 10299 2787 10308
rect 5092 10130 5120 11086
rect 5460 10810 5488 12718
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5538 12540 5846 12549
rect 5538 12538 5544 12540
rect 5600 12538 5624 12540
rect 5680 12538 5704 12540
rect 5760 12538 5784 12540
rect 5840 12538 5846 12540
rect 5600 12486 5602 12538
rect 5782 12486 5784 12538
rect 5538 12484 5544 12486
rect 5600 12484 5624 12486
rect 5680 12484 5704 12486
rect 5760 12484 5784 12486
rect 5840 12484 5846 12486
rect 5538 12475 5846 12484
rect 5920 12186 5948 12582
rect 5644 12170 5948 12186
rect 6012 12170 6040 12582
rect 5632 12164 5948 12170
rect 5684 12158 5948 12164
rect 6000 12164 6052 12170
rect 5632 12106 5684 12112
rect 6000 12106 6052 12112
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5538 11452 5846 11461
rect 5538 11450 5544 11452
rect 5600 11450 5624 11452
rect 5680 11450 5704 11452
rect 5760 11450 5784 11452
rect 5840 11450 5846 11452
rect 5600 11398 5602 11450
rect 5782 11398 5784 11450
rect 5538 11396 5544 11398
rect 5600 11396 5624 11398
rect 5680 11396 5704 11398
rect 5760 11396 5784 11398
rect 5840 11396 5846 11398
rect 5538 11387 5846 11396
rect 5920 10810 5948 11698
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9654 3188 9862
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2479 9276 2787 9285
rect 2479 9274 2485 9276
rect 2541 9274 2565 9276
rect 2621 9274 2645 9276
rect 2701 9274 2725 9276
rect 2781 9274 2787 9276
rect 2541 9222 2543 9274
rect 2723 9222 2725 9274
rect 2479 9220 2485 9222
rect 2541 9220 2565 9222
rect 2621 9220 2645 9222
rect 2701 9220 2725 9222
rect 2781 9220 2787 9222
rect 2479 9211 2787 9220
rect 3252 9042 3280 9318
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8634 1532 8774
rect 2976 8634 3004 8842
rect 3344 8634 3372 9998
rect 4008 9820 4316 9829
rect 4008 9818 4014 9820
rect 4070 9818 4094 9820
rect 4150 9818 4174 9820
rect 4230 9818 4254 9820
rect 4310 9818 4316 9820
rect 4070 9766 4072 9818
rect 4252 9766 4254 9818
rect 4008 9764 4014 9766
rect 4070 9764 4094 9766
rect 4150 9764 4174 9766
rect 4230 9764 4254 9766
rect 4310 9764 4316 9766
rect 4008 9755 4316 9764
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 3436 8974 3464 9318
rect 4356 8974 4384 9318
rect 5092 9042 5120 10066
rect 5460 9722 5488 10746
rect 6196 10674 6224 11154
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5538 10364 5846 10373
rect 5538 10362 5544 10364
rect 5600 10362 5624 10364
rect 5680 10362 5704 10364
rect 5760 10362 5784 10364
rect 5840 10362 5846 10364
rect 5600 10310 5602 10362
rect 5782 10310 5784 10362
rect 5538 10308 5544 10310
rect 5600 10308 5624 10310
rect 5680 10308 5704 10310
rect 5760 10308 5784 10310
rect 5840 10308 5846 10310
rect 5538 10299 5846 10308
rect 5920 10130 5948 10406
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9722 6040 9930
rect 5448 9716 5500 9722
rect 5276 9664 5448 9674
rect 5276 9658 5500 9664
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5276 9646 5488 9658
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 5778 1440 6802
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 2056 4078 2084 8570
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2412 8424 2464 8430
rect 2332 8372 2412 8378
rect 2332 8366 2464 8372
rect 2332 8350 2452 8366
rect 2332 7818 2360 8350
rect 2792 8294 2820 8434
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2479 8188 2787 8197
rect 2479 8186 2485 8188
rect 2541 8186 2565 8188
rect 2621 8186 2645 8188
rect 2701 8186 2725 8188
rect 2781 8186 2787 8188
rect 2541 8134 2543 8186
rect 2723 8134 2725 8186
rect 2479 8132 2485 8134
rect 2541 8132 2565 8134
rect 2621 8132 2645 8134
rect 2701 8132 2725 8134
rect 2781 8132 2787 8134
rect 2479 8123 2787 8132
rect 2884 8090 2912 8434
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 8016 2832 8022
rect 2976 7970 3004 8230
rect 2832 7964 3004 7970
rect 2780 7958 3004 7964
rect 2792 7942 3004 7958
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7002 2268 7686
rect 2332 7410 2360 7754
rect 2424 7546 2452 7822
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2792 7206 2820 7942
rect 3344 7886 3372 8434
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3160 7410 3188 7822
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2479 7100 2787 7109
rect 2479 7098 2485 7100
rect 2541 7098 2565 7100
rect 2621 7098 2645 7100
rect 2701 7098 2725 7100
rect 2781 7098 2787 7100
rect 2541 7046 2543 7098
rect 2723 7046 2725 7098
rect 2479 7044 2485 7046
rect 2541 7044 2565 7046
rect 2621 7044 2645 7046
rect 2701 7044 2725 7046
rect 2781 7044 2787 7046
rect 2479 7035 2787 7044
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 6322 3004 6734
rect 3160 6662 3188 7346
rect 3436 6798 3464 8910
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8498 3832 8842
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3804 8090 3832 8434
rect 3896 8362 3924 8774
rect 4008 8732 4316 8741
rect 4008 8730 4014 8732
rect 4070 8730 4094 8732
rect 4150 8730 4174 8732
rect 4230 8730 4254 8732
rect 4310 8730 4316 8732
rect 4070 8678 4072 8730
rect 4252 8678 4254 8730
rect 4008 8676 4014 8678
rect 4070 8676 4094 8678
rect 4150 8676 4174 8678
rect 4230 8676 4254 8678
rect 4310 8676 4316 8678
rect 4008 8667 4316 8676
rect 4356 8634 4384 8910
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4540 8514 4568 8774
rect 4356 8498 4568 8514
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4344 8492 4568 8498
rect 4396 8486 4568 8492
rect 4344 8434 4396 8440
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2148 5778 2176 6054
rect 2479 6012 2787 6021
rect 2479 6010 2485 6012
rect 2541 6010 2565 6012
rect 2621 6010 2645 6012
rect 2701 6010 2725 6012
rect 2781 6010 2787 6012
rect 2541 5958 2543 6010
rect 2723 5958 2725 6010
rect 2479 5956 2485 5958
rect 2541 5956 2565 5958
rect 2621 5956 2645 5958
rect 2701 5956 2725 5958
rect 2781 5956 2787 5958
rect 2479 5947 2787 5956
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2884 5710 2912 6054
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2976 5166 3004 6258
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5370 3096 6190
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4622 2176 4966
rect 2479 4924 2787 4933
rect 2479 4922 2485 4924
rect 2541 4922 2565 4924
rect 2621 4922 2645 4924
rect 2701 4922 2725 4924
rect 2781 4922 2787 4924
rect 2541 4870 2543 4922
rect 2723 4870 2725 4922
rect 2479 4868 2485 4870
rect 2541 4868 2565 4870
rect 2621 4868 2645 4870
rect 2701 4868 2725 4870
rect 2781 4868 2787 4870
rect 2479 4859 2787 4868
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2320 4140 2372 4146
rect 2240 4100 2320 4128
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2056 3602 2084 4014
rect 2240 3670 2268 4100
rect 2320 4082 2372 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2884 4026 2912 4082
rect 2884 3998 3096 4026
rect 3160 4010 3188 6598
rect 3712 6118 3740 6666
rect 3896 6322 3924 8298
rect 4356 7886 4384 8434
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4008 7644 4316 7653
rect 4008 7642 4014 7644
rect 4070 7642 4094 7644
rect 4150 7642 4174 7644
rect 4230 7642 4254 7644
rect 4310 7642 4316 7644
rect 4070 7590 4072 7642
rect 4252 7590 4254 7642
rect 4008 7588 4014 7590
rect 4070 7588 4094 7590
rect 4150 7588 4174 7590
rect 4230 7588 4254 7590
rect 4310 7588 4316 7590
rect 4008 7579 4316 7588
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4008 6556 4316 6565
rect 4008 6554 4014 6556
rect 4070 6554 4094 6556
rect 4150 6554 4174 6556
rect 4230 6554 4254 6556
rect 4310 6554 4316 6556
rect 4070 6502 4072 6554
rect 4252 6502 4254 6554
rect 4008 6500 4014 6502
rect 4070 6500 4094 6502
rect 4150 6500 4174 6502
rect 4230 6500 4254 6502
rect 4310 6500 4316 6502
rect 4008 6491 4316 6500
rect 4356 6390 4384 6666
rect 4448 6458 4476 6666
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3344 5234 3372 6054
rect 3804 5930 3832 6054
rect 3712 5902 3832 5930
rect 3712 5574 3740 5902
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 5234 3740 5510
rect 3896 5302 3924 6258
rect 4344 6248 4396 6254
rect 4264 6208 4344 6236
rect 4264 5914 4292 6208
rect 4344 6190 4396 6196
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5914 4384 6054
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4008 5468 4316 5477
rect 4008 5466 4014 5468
rect 4070 5466 4094 5468
rect 4150 5466 4174 5468
rect 4230 5466 4254 5468
rect 4310 5466 4316 5468
rect 4070 5414 4072 5466
rect 4252 5414 4254 5466
rect 4008 5412 4014 5414
rect 4070 5412 4094 5414
rect 4150 5412 4174 5414
rect 4230 5412 4254 5414
rect 4310 5412 4316 5414
rect 4008 5403 4316 5412
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3712 5114 3740 5170
rect 3712 5086 3832 5114
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3068 3942 3096 3998
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2479 3836 2787 3845
rect 2479 3834 2485 3836
rect 2541 3834 2565 3836
rect 2621 3834 2645 3836
rect 2701 3834 2725 3836
rect 2781 3834 2787 3836
rect 2541 3782 2543 3834
rect 2723 3782 2725 3834
rect 2479 3780 2485 3782
rect 2541 3780 2565 3782
rect 2621 3780 2645 3782
rect 2701 3780 2725 3782
rect 2781 3780 2787 3782
rect 2479 3771 2787 3780
rect 2884 3738 2912 3878
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2228 3664 2280 3670
rect 2228 3606 2280 3612
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1596 2650 1624 3538
rect 2056 3398 2084 3538
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2884 3194 2912 3334
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2976 3058 3004 3878
rect 3160 3602 3188 3946
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3670 3372 3878
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3620 3534 3648 4218
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3942 3740 4014
rect 3804 3942 3832 5086
rect 4356 5030 4384 5850
rect 4448 5778 4476 6394
rect 4540 5778 4568 6598
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4008 4380 4316 4389
rect 4008 4378 4014 4380
rect 4070 4378 4094 4380
rect 4150 4378 4174 4380
rect 4230 4378 4254 4380
rect 4310 4378 4316 4380
rect 4070 4326 4072 4378
rect 4252 4326 4254 4378
rect 4008 4324 4014 4326
rect 4070 4324 4094 4326
rect 4150 4324 4174 4326
rect 4230 4324 4254 4326
rect 4310 4324 4316 4326
rect 4008 4315 4316 4324
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4080 4010 4108 4150
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3068 3194 3096 3470
rect 3056 3188 3108 3194
rect 3108 3148 3464 3176
rect 3056 3130 3108 3136
rect 3436 3058 3464 3148
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 2479 2748 2787 2757
rect 2479 2746 2485 2748
rect 2541 2746 2565 2748
rect 2621 2746 2645 2748
rect 2701 2746 2725 2748
rect 2781 2746 2787 2748
rect 2541 2694 2543 2746
rect 2723 2694 2725 2746
rect 2479 2692 2485 2694
rect 2541 2692 2565 2694
rect 2621 2692 2645 2694
rect 2701 2692 2725 2694
rect 2781 2692 2787 2694
rect 2479 2683 2787 2692
rect 2884 2650 2912 2994
rect 3620 2774 3648 3470
rect 3712 2990 3740 3878
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3804 2922 3832 3878
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3896 3074 3924 3606
rect 4264 3534 4292 3946
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4008 3292 4316 3301
rect 4008 3290 4014 3292
rect 4070 3290 4094 3292
rect 4150 3290 4174 3292
rect 4230 3290 4254 3292
rect 4310 3290 4316 3292
rect 4070 3238 4072 3290
rect 4252 3238 4254 3290
rect 4008 3236 4014 3238
rect 4070 3236 4094 3238
rect 4150 3236 4174 3238
rect 4230 3236 4254 3238
rect 4310 3236 4316 3238
rect 4008 3227 4316 3236
rect 4356 3194 4384 3878
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4264 3074 4292 3130
rect 4632 3074 4660 8502
rect 5092 8090 5120 8978
rect 5184 8906 5212 8978
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8566 5212 8842
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5276 8412 5304 9646
rect 5538 9276 5846 9285
rect 5538 9274 5544 9276
rect 5600 9274 5624 9276
rect 5680 9274 5704 9276
rect 5760 9274 5784 9276
rect 5840 9274 5846 9276
rect 5600 9222 5602 9274
rect 5782 9222 5784 9274
rect 5538 9220 5544 9222
rect 5600 9220 5624 9222
rect 5680 9220 5704 9222
rect 5760 9220 5784 9222
rect 5840 9220 5846 9222
rect 5538 9211 5846 9220
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5184 8384 5304 8412
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6458 4752 6598
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4816 6118 4844 7142
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4908 5914 4936 6734
rect 5000 6458 5028 7210
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5370 5028 6394
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5184 5098 5212 8384
rect 5460 6866 5488 8910
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8634 5764 8842
rect 6104 8634 6132 8978
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5538 8188 5846 8197
rect 5538 8186 5544 8188
rect 5600 8186 5624 8188
rect 5680 8186 5704 8188
rect 5760 8186 5784 8188
rect 5840 8186 5846 8188
rect 5600 8134 5602 8186
rect 5782 8134 5784 8186
rect 5538 8132 5544 8134
rect 5600 8132 5624 8134
rect 5680 8132 5704 8134
rect 5760 8132 5784 8134
rect 5840 8132 5846 8134
rect 5538 8123 5846 8132
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 5828 7262 5948 7290
rect 5828 7206 5856 7262
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5538 7100 5846 7109
rect 5538 7098 5544 7100
rect 5600 7098 5624 7100
rect 5680 7098 5704 7100
rect 5760 7098 5784 7100
rect 5840 7098 5846 7100
rect 5600 7046 5602 7098
rect 5782 7046 5784 7098
rect 5538 7044 5544 7046
rect 5600 7044 5624 7046
rect 5680 7044 5704 7046
rect 5760 7044 5784 7046
rect 5840 7044 5846 7046
rect 5538 7035 5846 7044
rect 5920 7002 5948 7262
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5908 6860 5960 6866
rect 6012 6848 6040 7142
rect 5960 6820 6040 6848
rect 5908 6802 5960 6808
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5370 5304 6190
rect 5368 5522 5396 6666
rect 5460 5846 5488 6802
rect 6104 6730 6132 7414
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5538 6012 5846 6021
rect 5538 6010 5544 6012
rect 5600 6010 5624 6012
rect 5680 6010 5704 6012
rect 5760 6010 5784 6012
rect 5840 6010 5846 6012
rect 5600 5958 5602 6010
rect 5782 5958 5784 6010
rect 5538 5956 5544 5958
rect 5600 5956 5624 5958
rect 5680 5956 5704 5958
rect 5760 5956 5784 5958
rect 5840 5956 5846 5958
rect 5538 5947 5846 5956
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5368 5494 5580 5522
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 4690 5212 5034
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4724 3126 4752 3946
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4908 3194 4936 4082
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5000 3126 5028 4082
rect 5276 4010 5304 5306
rect 5552 5302 5580 5494
rect 5920 5370 5948 6326
rect 6196 6118 6224 7210
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5534 6224 6054
rect 6288 5914 6316 13874
rect 8597 13628 8905 13637
rect 8597 13626 8603 13628
rect 8659 13626 8683 13628
rect 8739 13626 8763 13628
rect 8819 13626 8843 13628
rect 8899 13626 8905 13628
rect 8659 13574 8661 13626
rect 8841 13574 8843 13626
rect 8597 13572 8603 13574
rect 8659 13572 8683 13574
rect 8739 13572 8763 13574
rect 8819 13572 8843 13574
rect 8899 13572 8905 13574
rect 8597 13563 8905 13572
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 12918 6776 13330
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 6932 12918 6960 13262
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7067 13084 7375 13093
rect 7067 13082 7073 13084
rect 7129 13082 7153 13084
rect 7209 13082 7233 13084
rect 7289 13082 7313 13084
rect 7369 13082 7375 13084
rect 7129 13030 7131 13082
rect 7311 13030 7313 13082
rect 7067 13028 7073 13030
rect 7129 13028 7153 13030
rect 7209 13028 7233 13030
rect 7289 13028 7313 13030
rect 7369 13028 7375 13030
rect 7067 13019 7375 13028
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 8566 6408 12038
rect 6564 11898 6592 12582
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6656 11354 6684 12854
rect 6748 12170 6776 12854
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10742 6684 10950
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6748 10538 6776 12106
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11694 6868 12038
rect 6932 11694 6960 12854
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12442 7328 12786
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7300 12186 7328 12378
rect 7392 12306 7420 12582
rect 7484 12442 7512 13126
rect 7760 12782 7788 13126
rect 7852 12918 7880 13126
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 8128 12442 8156 13262
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8022 12336 8078 12345
rect 7380 12300 7432 12306
rect 8220 12306 8248 12582
rect 8496 12442 8524 12854
rect 8597 12540 8905 12549
rect 8597 12538 8603 12540
rect 8659 12538 8683 12540
rect 8739 12538 8763 12540
rect 8819 12538 8843 12540
rect 8899 12538 8905 12540
rect 8659 12486 8661 12538
rect 8841 12486 8843 12538
rect 8597 12484 8603 12486
rect 8659 12484 8683 12486
rect 8739 12484 8763 12486
rect 8819 12484 8843 12486
rect 8899 12484 8905 12486
rect 8597 12475 8905 12484
rect 9140 12442 9168 13262
rect 9784 12986 9812 13262
rect 10126 13084 10434 13093
rect 10126 13082 10132 13084
rect 10188 13082 10212 13084
rect 10268 13082 10292 13084
rect 10348 13082 10372 13084
rect 10428 13082 10434 13084
rect 10188 13030 10190 13082
rect 10370 13030 10372 13082
rect 10126 13028 10132 13030
rect 10188 13028 10212 13030
rect 10268 13028 10292 13030
rect 10348 13028 10372 13030
rect 10428 13028 10434 13030
rect 10126 13019 10434 13028
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 9784 12442 9812 12786
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 8022 12271 8078 12280
rect 8208 12300 8260 12306
rect 7380 12242 7432 12248
rect 8036 12238 8064 12271
rect 8208 12242 8260 12248
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 8024 12232 8076 12238
rect 7300 12158 7512 12186
rect 8024 12174 8076 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 7067 11996 7375 12005
rect 7067 11994 7073 11996
rect 7129 11994 7153 11996
rect 7209 11994 7233 11996
rect 7289 11994 7313 11996
rect 7369 11994 7375 11996
rect 7129 11942 7131 11994
rect 7311 11942 7313 11994
rect 7067 11940 7073 11942
rect 7129 11940 7153 11942
rect 7209 11940 7233 11942
rect 7289 11940 7313 11942
rect 7369 11940 7375 11942
rect 7067 11931 7375 11940
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6840 11370 6868 11630
rect 6840 11354 6960 11370
rect 6840 11348 6972 11354
rect 6840 11342 6920 11348
rect 6920 11290 6972 11296
rect 7024 11286 7052 11698
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7208 11218 7236 11494
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10792 6960 11086
rect 7208 11014 7236 11154
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7067 10908 7375 10917
rect 7067 10906 7073 10908
rect 7129 10906 7153 10908
rect 7209 10906 7233 10908
rect 7289 10906 7313 10908
rect 7369 10906 7375 10908
rect 7129 10854 7131 10906
rect 7311 10854 7313 10906
rect 7067 10852 7073 10854
rect 7129 10852 7153 10854
rect 7209 10852 7233 10854
rect 7289 10852 7313 10854
rect 7369 10852 7375 10854
rect 7067 10843 7375 10852
rect 6932 10764 7144 10792
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 7024 10266 7052 10610
rect 7116 10606 7144 10764
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7116 10130 7144 10542
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7067 9820 7375 9829
rect 7067 9818 7073 9820
rect 7129 9818 7153 9820
rect 7209 9818 7233 9820
rect 7289 9818 7313 9820
rect 7369 9818 7375 9820
rect 7129 9766 7131 9818
rect 7311 9766 7313 9818
rect 7067 9764 7073 9766
rect 7129 9764 7153 9766
rect 7209 9764 7233 9766
rect 7289 9764 7313 9766
rect 7369 9764 7375 9766
rect 7067 9755 7375 9764
rect 7484 9722 7512 12158
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11354 7604 12038
rect 9140 11898 9168 12174
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7760 10674 7788 11086
rect 8036 11082 8064 11494
rect 8597 11452 8905 11461
rect 8597 11450 8603 11452
rect 8659 11450 8683 11452
rect 8739 11450 8763 11452
rect 8819 11450 8843 11452
rect 8899 11450 8905 11452
rect 8659 11398 8661 11450
rect 8841 11398 8843 11450
rect 8597 11396 8603 11398
rect 8659 11396 8683 11398
rect 8739 11396 8763 11398
rect 8819 11396 8843 11398
rect 8899 11396 8905 11398
rect 8597 11387 8905 11396
rect 9324 11354 9352 12106
rect 9508 11694 9536 12174
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11150 9444 11494
rect 9600 11234 9628 11698
rect 9508 11206 9628 11234
rect 9508 11150 9536 11206
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8036 10674 8064 11018
rect 8404 10742 8432 11018
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7760 9926 7788 10610
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8974 7420 9318
rect 7576 8974 7604 9522
rect 7760 9178 7788 9862
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7067 8732 7375 8741
rect 7067 8730 7073 8732
rect 7129 8730 7153 8732
rect 7209 8730 7233 8732
rect 7289 8730 7313 8732
rect 7369 8730 7375 8732
rect 7129 8678 7131 8730
rect 7311 8678 7313 8730
rect 7067 8676 7073 8678
rect 7129 8676 7153 8678
rect 7209 8676 7233 8678
rect 7289 8676 7313 8678
rect 7369 8676 7375 8678
rect 7067 8667 7375 8676
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7886 7696 8230
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6730 6592 7142
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6656 5710 6684 7822
rect 7067 7644 7375 7653
rect 7067 7642 7073 7644
rect 7129 7642 7153 7644
rect 7209 7642 7233 7644
rect 7289 7642 7313 7644
rect 7369 7642 7375 7644
rect 7129 7590 7131 7642
rect 7311 7590 7313 7642
rect 7067 7588 7073 7590
rect 7129 7588 7153 7590
rect 7209 7588 7233 7590
rect 7289 7588 7313 7590
rect 7369 7588 7375 7590
rect 7067 7579 7375 7588
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6798 7604 7142
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7067 6556 7375 6565
rect 7067 6554 7073 6556
rect 7129 6554 7153 6556
rect 7209 6554 7233 6556
rect 7289 6554 7313 6556
rect 7369 6554 7375 6556
rect 7129 6502 7131 6554
rect 7311 6502 7313 6554
rect 7067 6500 7073 6502
rect 7129 6500 7153 6502
rect 7209 6500 7233 6502
rect 7289 6500 7313 6502
rect 7369 6500 7375 6502
rect 7067 6491 7375 6500
rect 7576 6390 7604 6734
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6104 5506 6224 5534
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 6104 5234 6132 5506
rect 7067 5468 7375 5477
rect 7067 5466 7073 5468
rect 7129 5466 7153 5468
rect 7209 5466 7233 5468
rect 7289 5466 7313 5468
rect 7369 5466 7375 5468
rect 7129 5414 7131 5466
rect 7311 5414 7313 5466
rect 7067 5412 7073 5414
rect 7129 5412 7153 5414
rect 7209 5412 7233 5414
rect 7289 5412 7313 5414
rect 7369 5412 7375 5414
rect 7067 5403 7375 5412
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5538 4924 5846 4933
rect 5538 4922 5544 4924
rect 5600 4922 5624 4924
rect 5680 4922 5704 4924
rect 5760 4922 5784 4924
rect 5840 4922 5846 4924
rect 5600 4870 5602 4922
rect 5782 4870 5784 4922
rect 5538 4868 5544 4870
rect 5600 4868 5624 4870
rect 5680 4868 5704 4870
rect 5760 4868 5784 4870
rect 5840 4868 5846 4870
rect 5538 4859 5846 4868
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6932 4128 6960 5238
rect 7484 5234 7512 5850
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7067 4380 7375 4389
rect 7067 4378 7073 4380
rect 7129 4378 7153 4380
rect 7209 4378 7233 4380
rect 7289 4378 7313 4380
rect 7369 4378 7375 4380
rect 7129 4326 7131 4378
rect 7311 4326 7313 4378
rect 7067 4324 7073 4326
rect 7129 4324 7153 4326
rect 7209 4324 7233 4326
rect 7289 4324 7313 4326
rect 7369 4324 7375 4326
rect 7067 4315 7375 4324
rect 7288 4140 7340 4146
rect 6932 4100 7288 4128
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5276 3534 5304 3946
rect 5538 3836 5846 3845
rect 5538 3834 5544 3836
rect 5600 3834 5624 3836
rect 5680 3834 5704 3836
rect 5760 3834 5784 3836
rect 5840 3834 5846 3836
rect 5600 3782 5602 3834
rect 5782 3782 5784 3834
rect 5538 3780 5544 3782
rect 5600 3780 5624 3782
rect 5680 3780 5704 3782
rect 5760 3780 5784 3782
rect 5840 3780 5846 3782
rect 5538 3771 5846 3780
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5080 3528 5132 3534
rect 5264 3528 5316 3534
rect 5080 3470 5132 3476
rect 5184 3488 5264 3516
rect 3896 3058 4016 3074
rect 3896 3052 4028 3058
rect 3896 3046 3976 3052
rect 4264 3046 4660 3074
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 3976 2994 4028 3000
rect 4632 2990 4660 3046
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 3620 2746 3740 2774
rect 3712 2650 3740 2746
rect 4356 2650 4384 2858
rect 4908 2650 4936 2926
rect 5092 2922 5120 3470
rect 5184 3058 5212 3488
rect 5264 3470 5316 3476
rect 5460 3194 5488 3606
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5920 3194 5948 4014
rect 6012 3602 6040 4014
rect 6104 3670 6132 4082
rect 6644 4072 6696 4078
rect 6642 4040 6644 4049
rect 6828 4072 6880 4078
rect 6696 4040 6698 4049
rect 6828 4014 6880 4020
rect 6642 3975 6698 3984
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6104 3074 6132 3606
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 3194 6316 3538
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6184 3120 6236 3126
rect 6104 3068 6184 3074
rect 6104 3062 6236 3068
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 6104 3046 6224 3062
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5538 2748 5846 2757
rect 5538 2746 5544 2748
rect 5600 2746 5624 2748
rect 5680 2746 5704 2748
rect 5760 2746 5784 2748
rect 5840 2746 5846 2748
rect 5600 2694 5602 2746
rect 5782 2694 5784 2746
rect 5538 2692 5544 2694
rect 5600 2692 5624 2694
rect 5680 2692 5704 2694
rect 5760 2692 5784 2694
rect 5840 2692 5846 2694
rect 5538 2683 5846 2692
rect 6104 2650 6132 3046
rect 6288 2922 6316 3130
rect 6380 3058 6408 3470
rect 6656 3194 6684 3878
rect 6748 3602 6776 3878
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3602 6960 4100
rect 7576 4128 7604 6326
rect 7760 5534 7788 9114
rect 8036 8498 8064 10610
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 9722 8248 10406
rect 8597 10364 8905 10373
rect 8597 10362 8603 10364
rect 8659 10362 8683 10364
rect 8739 10362 8763 10364
rect 8819 10362 8843 10364
rect 8899 10362 8905 10364
rect 8659 10310 8661 10362
rect 8841 10310 8843 10362
rect 8597 10308 8603 10310
rect 8659 10308 8683 10310
rect 8739 10308 8763 10310
rect 8819 10308 8843 10310
rect 8899 10308 8905 10310
rect 8597 10299 8905 10308
rect 9416 10266 9444 11086
rect 9508 10810 9536 11086
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9692 10742 9720 12242
rect 9876 12170 9904 12718
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12374 10088 12650
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12374 10180 12582
rect 10796 12442 10824 12786
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10140 12368 10192 12374
rect 10232 12368 10284 12374
rect 10140 12310 10192 12316
rect 10230 12336 10232 12345
rect 10284 12336 10286 12345
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11778 9996 12038
rect 10060 11898 10088 12310
rect 10230 12271 10286 12280
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10126 11996 10434 12005
rect 10126 11994 10132 11996
rect 10188 11994 10212 11996
rect 10268 11994 10292 11996
rect 10348 11994 10372 11996
rect 10428 11994 10434 11996
rect 10188 11942 10190 11994
rect 10370 11942 10372 11994
rect 10126 11940 10132 11942
rect 10188 11940 10212 11942
rect 10268 11940 10292 11942
rect 10348 11940 10372 11942
rect 10428 11940 10434 11942
rect 10126 11931 10434 11940
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9968 11762 10180 11778
rect 10520 11762 10548 12038
rect 9968 11756 10192 11762
rect 9968 11750 10140 11756
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9784 11218 9812 11562
rect 9968 11354 9996 11750
rect 10140 11698 10192 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10336 11642 10364 11698
rect 10244 11614 10364 11642
rect 10244 11558 10272 11614
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 10060 10674 10088 10950
rect 10126 10908 10434 10917
rect 10126 10906 10132 10908
rect 10188 10906 10212 10908
rect 10268 10906 10292 10908
rect 10348 10906 10372 10908
rect 10428 10906 10434 10908
rect 10188 10854 10190 10906
rect 10370 10854 10372 10906
rect 10126 10852 10132 10854
rect 10188 10852 10212 10854
rect 10268 10852 10292 10854
rect 10348 10852 10372 10854
rect 10428 10852 10434 10854
rect 10126 10843 10434 10852
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9784 10266 9812 10610
rect 10140 10600 10192 10606
rect 10060 10548 10140 10554
rect 10060 10542 10192 10548
rect 10060 10526 10180 10542
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8496 9178 8524 9590
rect 9784 9586 9812 10202
rect 10060 9994 10088 10526
rect 10520 10266 10548 11086
rect 10704 10810 10732 11494
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 10266 10640 10474
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9968 9518 9996 9862
rect 10060 9586 10088 9930
rect 10126 9820 10434 9829
rect 10126 9818 10132 9820
rect 10188 9818 10212 9820
rect 10268 9818 10292 9820
rect 10348 9818 10372 9820
rect 10428 9818 10434 9820
rect 10188 9766 10190 9818
rect 10370 9766 10372 9818
rect 10126 9764 10132 9766
rect 10188 9764 10212 9766
rect 10268 9764 10292 9766
rect 10348 9764 10372 9766
rect 10428 9764 10434 9766
rect 10126 9755 10434 9764
rect 10520 9654 10548 10202
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10704 9382 10732 9522
rect 10888 9450 10916 11154
rect 10980 9586 11008 13874
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 11656 13628 11964 13637
rect 11656 13626 11662 13628
rect 11718 13626 11742 13628
rect 11798 13626 11822 13628
rect 11878 13626 11902 13628
rect 11958 13626 11964 13628
rect 11718 13574 11720 13626
rect 11900 13574 11902 13626
rect 11656 13572 11662 13574
rect 11718 13572 11742 13574
rect 11798 13572 11822 13574
rect 11878 13572 11902 13574
rect 11958 13572 11964 13574
rect 11656 13563 11964 13572
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11656 12540 11964 12549
rect 11656 12538 11662 12540
rect 11718 12538 11742 12540
rect 11798 12538 11822 12540
rect 11878 12538 11902 12540
rect 11958 12538 11964 12540
rect 11718 12486 11720 12538
rect 11900 12486 11902 12538
rect 11656 12484 11662 12486
rect 11718 12484 11742 12486
rect 11798 12484 11822 12486
rect 11878 12484 11902 12486
rect 11958 12484 11964 12486
rect 11656 12475 11964 12484
rect 11992 12442 12020 13126
rect 12728 12918 12756 13738
rect 13185 13084 13493 13093
rect 13185 13082 13191 13084
rect 13247 13082 13271 13084
rect 13327 13082 13351 13084
rect 13407 13082 13431 13084
rect 13487 13082 13493 13084
rect 13247 13030 13249 13082
rect 13429 13030 13431 13082
rect 13185 13028 13191 13030
rect 13247 13028 13271 13030
rect 13327 13028 13351 13030
rect 13407 13028 13431 13030
rect 13487 13028 13493 13030
rect 13185 13019 13493 13028
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11164 11354 11192 11630
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11072 10606 11100 11290
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11164 10810 11192 11018
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11164 9654 11192 10746
rect 11256 10062 11284 11494
rect 11348 11150 11376 11494
rect 11440 11354 11468 12174
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11694 11560 12038
rect 11992 11898 12020 12378
rect 12728 12306 12756 12854
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 13185 11996 13493 12005
rect 13185 11994 13191 11996
rect 13247 11994 13271 11996
rect 13327 11994 13351 11996
rect 13407 11994 13431 11996
rect 13487 11994 13493 11996
rect 13247 11942 13249 11994
rect 13429 11942 13431 11994
rect 13185 11940 13191 11942
rect 13247 11940 13271 11942
rect 13327 11940 13351 11942
rect 13407 11940 13431 11942
rect 13487 11940 13493 11942
rect 13185 11931 13493 11940
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11532 11150 11560 11630
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11656 11452 11964 11461
rect 11656 11450 11662 11452
rect 11718 11450 11742 11452
rect 11798 11450 11822 11452
rect 11878 11450 11902 11452
rect 11958 11450 11964 11452
rect 11718 11398 11720 11450
rect 11900 11398 11902 11450
rect 11656 11396 11662 11398
rect 11718 11396 11742 11398
rect 11798 11396 11822 11398
rect 11878 11396 11902 11398
rect 11958 11396 11964 11398
rect 11656 11387 11964 11396
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 11054 11652 11086
rect 11624 11026 11836 11054
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10674 11560 10950
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11808 10538 11836 11026
rect 11992 10810 12020 11494
rect 12268 11150 12296 11494
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11980 10804 12032 10810
rect 12032 10764 12112 10792
rect 11980 10746 12032 10752
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11440 9586 11468 10406
rect 11532 10266 11560 10474
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11656 10364 11964 10373
rect 11656 10362 11662 10364
rect 11718 10362 11742 10364
rect 11798 10362 11822 10364
rect 11878 10362 11902 10364
rect 11958 10362 11964 10364
rect 11718 10310 11720 10362
rect 11900 10310 11902 10362
rect 11656 10308 11662 10310
rect 11718 10308 11742 10310
rect 11798 10308 11822 10310
rect 11878 10308 11902 10310
rect 11958 10308 11964 10310
rect 11656 10299 11964 10308
rect 11992 10266 12020 10406
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12084 10062 12112 10764
rect 12176 10266 12204 11086
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12268 10062 12296 10474
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9602 11652 9658
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11532 9574 11652 9602
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 8597 9276 8905 9285
rect 8597 9274 8603 9276
rect 8659 9274 8683 9276
rect 8739 9274 8763 9276
rect 8819 9274 8843 9276
rect 8899 9274 8905 9276
rect 8659 9222 8661 9274
rect 8841 9222 8843 9274
rect 8597 9220 8603 9222
rect 8659 9220 8683 9222
rect 8739 9220 8763 9222
rect 8819 9220 8843 9222
rect 8899 9220 8905 9222
rect 8597 9211 8905 9220
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7668 5506 7788 5534
rect 8220 5534 8248 8434
rect 8312 7750 8340 8774
rect 10126 8732 10434 8741
rect 10126 8730 10132 8732
rect 10188 8730 10212 8732
rect 10268 8730 10292 8732
rect 10348 8730 10372 8732
rect 10428 8730 10434 8732
rect 10188 8678 10190 8730
rect 10370 8678 10372 8730
rect 10126 8676 10132 8678
rect 10188 8676 10212 8678
rect 10268 8676 10292 8678
rect 10348 8676 10372 8678
rect 10428 8676 10434 8678
rect 10126 8667 10434 8676
rect 10520 8498 10548 9318
rect 11532 9110 11560 9574
rect 11656 9276 11964 9285
rect 11656 9274 11662 9276
rect 11718 9274 11742 9276
rect 11798 9274 11822 9276
rect 11878 9274 11902 9276
rect 11958 9274 11964 9276
rect 11718 9222 11720 9274
rect 11900 9222 11902 9274
rect 11656 9220 11662 9222
rect 11718 9220 11742 9222
rect 11798 9220 11822 9222
rect 11878 9220 11902 9222
rect 11958 9220 11964 9222
rect 11656 9211 11964 9220
rect 12360 9178 12388 11086
rect 13185 10908 13493 10917
rect 13185 10906 13191 10908
rect 13247 10906 13271 10908
rect 13327 10906 13351 10908
rect 13407 10906 13431 10908
rect 13487 10906 13493 10908
rect 13247 10854 13249 10906
rect 13429 10854 13431 10906
rect 13185 10852 13191 10854
rect 13247 10852 13271 10854
rect 13327 10852 13351 10854
rect 13407 10852 13431 10854
rect 13487 10852 13493 10854
rect 13185 10843 13493 10852
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12636 10062 12664 10542
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12728 9586 12756 10202
rect 13004 10169 13032 10542
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 13185 9820 13493 9829
rect 13185 9818 13191 9820
rect 13247 9818 13271 9820
rect 13327 9818 13351 9820
rect 13407 9818 13431 9820
rect 13487 9818 13493 9820
rect 13247 9766 13249 9818
rect 13429 9766 13431 9818
rect 13185 9764 13191 9766
rect 13247 9764 13271 9766
rect 13327 9764 13351 9766
rect 13407 9764 13431 9766
rect 13487 9764 13493 9766
rect 13185 9755 13493 9764
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 8597 8188 8905 8197
rect 8597 8186 8603 8188
rect 8659 8186 8683 8188
rect 8739 8186 8763 8188
rect 8819 8186 8843 8188
rect 8899 8186 8905 8188
rect 8659 8134 8661 8186
rect 8841 8134 8843 8186
rect 8597 8132 8603 8134
rect 8659 8132 8683 8134
rect 8739 8132 8763 8134
rect 8819 8132 8843 8134
rect 8899 8132 8905 8134
rect 8597 8123 8905 8132
rect 11440 7954 11468 8774
rect 12360 8634 12388 8910
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11656 8188 11964 8197
rect 11656 8186 11662 8188
rect 11718 8186 11742 8188
rect 11798 8186 11822 8188
rect 11878 8186 11902 8188
rect 11958 8186 11964 8188
rect 11718 8134 11720 8186
rect 11900 8134 11902 8186
rect 11656 8132 11662 8134
rect 11718 8132 11742 8134
rect 11798 8132 11822 8134
rect 11878 8132 11902 8134
rect 11958 8132 11964 8134
rect 11656 8123 11964 8132
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8312 6118 8340 7686
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7002 8524 7822
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8597 7100 8905 7109
rect 8597 7098 8603 7100
rect 8659 7098 8683 7100
rect 8739 7098 8763 7100
rect 8819 7098 8843 7100
rect 8899 7098 8905 7100
rect 8659 7046 8661 7098
rect 8841 7046 8843 7098
rect 8597 7044 8603 7046
rect 8659 7044 8683 7046
rect 8739 7044 8763 7046
rect 8819 7044 8843 7046
rect 8899 7044 8905 7046
rect 8597 7035 8905 7044
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8956 6798 8984 7754
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6798 9076 7346
rect 9232 7002 9260 7822
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6458 8432 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5710 8340 6054
rect 8597 6012 8905 6021
rect 8597 6010 8603 6012
rect 8659 6010 8683 6012
rect 8739 6010 8763 6012
rect 8819 6010 8843 6012
rect 8899 6010 8905 6012
rect 8659 5958 8661 6010
rect 8841 5958 8843 6010
rect 8597 5956 8603 5958
rect 8659 5956 8683 5958
rect 8739 5956 8763 5958
rect 8819 5956 8843 5958
rect 8899 5956 8905 5958
rect 8597 5947 8905 5956
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8220 5506 8340 5534
rect 7668 4282 7696 5506
rect 8312 5302 8340 5506
rect 8772 5370 8800 5850
rect 9048 5778 9076 6734
rect 9324 6730 9352 7686
rect 9416 7290 9444 7754
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 10126 7644 10434 7653
rect 10126 7642 10132 7644
rect 10188 7642 10212 7644
rect 10268 7642 10292 7644
rect 10348 7642 10372 7644
rect 10428 7642 10434 7644
rect 10188 7590 10190 7642
rect 10370 7590 10372 7642
rect 10126 7588 10132 7590
rect 10188 7588 10212 7590
rect 10268 7588 10292 7590
rect 10348 7588 10372 7590
rect 10428 7588 10434 7590
rect 10126 7579 10434 7588
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9416 7262 9536 7290
rect 9508 7206 9536 7262
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9508 6458 9536 7142
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9508 5370 9536 6394
rect 9600 6322 9628 6938
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9784 6458 9812 6734
rect 9876 6458 9904 6734
rect 10152 6730 10180 7142
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5370 9812 6190
rect 9876 5370 9904 6394
rect 10060 6322 10088 6598
rect 10126 6556 10434 6565
rect 10126 6554 10132 6556
rect 10188 6554 10212 6556
rect 10268 6554 10292 6556
rect 10348 6554 10372 6556
rect 10428 6554 10434 6556
rect 10188 6502 10190 6554
rect 10370 6502 10372 6554
rect 10126 6500 10132 6502
rect 10188 6500 10212 6502
rect 10268 6500 10292 6502
rect 10348 6500 10372 6502
rect 10428 6500 10434 6502
rect 10126 6491 10434 6500
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10126 5468 10434 5477
rect 10126 5466 10132 5468
rect 10188 5466 10212 5468
rect 10268 5466 10292 5468
rect 10348 5466 10372 5468
rect 10428 5466 10434 5468
rect 10188 5414 10190 5466
rect 10370 5414 10372 5466
rect 10126 5412 10132 5414
rect 10188 5412 10212 5414
rect 10268 5412 10292 5414
rect 10348 5412 10372 5414
rect 10428 5412 10434 5414
rect 10126 5403 10434 5412
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4282 8524 5170
rect 8597 4924 8905 4933
rect 8597 4922 8603 4924
rect 8659 4922 8683 4924
rect 8739 4922 8763 4924
rect 8819 4922 8843 4924
rect 8899 4922 8905 4924
rect 8659 4870 8661 4922
rect 8841 4870 8843 4922
rect 8597 4868 8603 4870
rect 8659 4868 8683 4870
rect 8739 4868 8763 4870
rect 8819 4868 8843 4870
rect 8899 4868 8905 4870
rect 8597 4859 8905 4868
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 9140 4214 9168 5238
rect 10796 5234 10824 6938
rect 11164 6866 11192 7822
rect 12176 7818 12204 8230
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12268 7342 12296 8434
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 11656 7100 11964 7109
rect 11656 7098 11662 7100
rect 11718 7098 11742 7100
rect 11798 7098 11822 7100
rect 11878 7098 11902 7100
rect 11958 7098 11964 7100
rect 11718 7046 11720 7098
rect 11900 7046 11902 7098
rect 11656 7044 11662 7046
rect 11718 7044 11742 7046
rect 11798 7044 11822 7046
rect 11878 7044 11902 7046
rect 11958 7044 11964 7046
rect 11656 7035 11964 7044
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 9232 4826 9260 5170
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 7656 4140 7708 4146
rect 7576 4100 7656 4128
rect 7288 4082 7340 4088
rect 7656 4082 7708 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7116 3738 7144 3946
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7024 3505 7052 3674
rect 7194 3632 7250 3641
rect 7116 3602 7194 3618
rect 7104 3596 7194 3602
rect 7156 3590 7194 3596
rect 7194 3567 7250 3576
rect 7104 3538 7156 3544
rect 7300 3534 7328 4082
rect 7668 4010 7696 4082
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7760 3670 7788 4082
rect 8036 3738 8064 4082
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7288 3528 7340 3534
rect 7010 3496 7066 3505
rect 6920 3460 6972 3466
rect 7288 3470 7340 3476
rect 7010 3431 7066 3440
rect 6920 3402 6972 3408
rect 6932 3194 6960 3402
rect 7760 3398 7788 3606
rect 7852 3505 7880 3606
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7838 3496 7894 3505
rect 7838 3431 7894 3440
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7067 3292 7375 3301
rect 7067 3290 7073 3292
rect 7129 3290 7153 3292
rect 7209 3290 7233 3292
rect 7289 3290 7313 3292
rect 7369 3290 7375 3292
rect 7129 3238 7131 3290
rect 7311 3238 7313 3290
rect 7067 3236 7073 3238
rect 7129 3236 7153 3238
rect 7209 3236 7233 3238
rect 7289 3236 7313 3238
rect 7369 3236 7375 3238
rect 7067 3227 7375 3236
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7484 3058 7512 3334
rect 7760 3194 7788 3334
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 2774 6316 2858
rect 6196 2746 6316 2774
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6196 2446 6224 2746
rect 6472 2650 6500 2994
rect 8036 2990 8064 3538
rect 8128 3194 8156 4082
rect 8404 3641 8432 4082
rect 9048 4026 9076 4082
rect 9140 4049 9168 4150
rect 8772 3998 9076 4026
rect 9126 4040 9182 4049
rect 8772 3942 8800 3998
rect 9126 3975 9182 3984
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 8597 3836 8905 3845
rect 8597 3834 8603 3836
rect 8659 3834 8683 3836
rect 8739 3834 8763 3836
rect 8819 3834 8843 3836
rect 8899 3834 8905 3836
rect 8659 3782 8661 3834
rect 8841 3782 8843 3834
rect 8597 3780 8603 3782
rect 8659 3780 8683 3782
rect 8739 3780 8763 3782
rect 8819 3780 8843 3782
rect 8899 3780 8905 3782
rect 8597 3771 8905 3780
rect 8390 3632 8446 3641
rect 8956 3602 8984 3878
rect 9048 3641 9076 3878
rect 9034 3632 9090 3641
rect 8390 3567 8446 3576
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8944 3596 8996 3602
rect 9034 3567 9036 3576
rect 8944 3538 8996 3544
rect 9088 3567 9090 3576
rect 9036 3538 9088 3544
rect 8482 3496 8538 3505
rect 8538 3466 8616 3482
rect 8538 3460 8628 3466
rect 8538 3454 8576 3460
rect 8482 3431 8538 3440
rect 8576 3402 8628 3408
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8220 3194 8248 3334
rect 8312 3194 8340 3334
rect 8588 3194 8616 3402
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8680 3126 8708 3538
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8864 2990 8892 3402
rect 9140 3194 9168 3878
rect 9324 3738 9352 3878
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3534 9444 4966
rect 9784 4146 9812 4966
rect 10704 4622 10732 5170
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10126 4380 10434 4389
rect 10126 4378 10132 4380
rect 10188 4378 10212 4380
rect 10268 4378 10292 4380
rect 10348 4378 10372 4380
rect 10428 4378 10434 4380
rect 10188 4326 10190 4378
rect 10370 4326 10372 4378
rect 10126 4324 10132 4326
rect 10188 4324 10212 4326
rect 10268 4324 10292 4326
rect 10348 4324 10372 4326
rect 10428 4324 10434 4326
rect 10126 4315 10434 4324
rect 10796 4282 10824 5170
rect 11164 4622 11192 6802
rect 12176 6730 12204 7142
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 11656 6012 11964 6021
rect 11656 6010 11662 6012
rect 11718 6010 11742 6012
rect 11798 6010 11822 6012
rect 11878 6010 11902 6012
rect 11958 6010 11964 6012
rect 11718 5958 11720 6010
rect 11900 5958 11902 6010
rect 11656 5956 11662 5958
rect 11718 5956 11742 5958
rect 11798 5956 11822 5958
rect 11878 5956 11902 5958
rect 11958 5956 11964 5958
rect 11656 5947 11964 5956
rect 12268 5534 12296 7278
rect 12176 5506 12296 5534
rect 12636 5534 12664 9318
rect 12728 6322 12756 9522
rect 13185 8732 13493 8741
rect 13185 8730 13191 8732
rect 13247 8730 13271 8732
rect 13327 8730 13351 8732
rect 13407 8730 13431 8732
rect 13487 8730 13493 8732
rect 13247 8678 13249 8730
rect 13429 8678 13431 8730
rect 13185 8676 13191 8678
rect 13247 8676 13271 8678
rect 13327 8676 13351 8678
rect 13407 8676 13431 8678
rect 13487 8676 13493 8678
rect 13185 8667 13493 8676
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 8090 12940 8366
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13185 7644 13493 7653
rect 13185 7642 13191 7644
rect 13247 7642 13271 7644
rect 13327 7642 13351 7644
rect 13407 7642 13431 7644
rect 13487 7642 13493 7644
rect 13247 7590 13249 7642
rect 13429 7590 13431 7642
rect 13185 7588 13191 7590
rect 13247 7588 13271 7590
rect 13327 7588 13351 7590
rect 13407 7588 13431 7590
rect 13487 7588 13493 7590
rect 13185 7579 13493 7588
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6390 12940 6598
rect 13185 6556 13493 6565
rect 13185 6554 13191 6556
rect 13247 6554 13271 6556
rect 13327 6554 13351 6556
rect 13407 6554 13431 6556
rect 13487 6554 13493 6556
rect 13247 6502 13249 6554
rect 13429 6502 13431 6554
rect 13185 6500 13191 6502
rect 13247 6500 13271 6502
rect 13327 6500 13351 6502
rect 13407 6500 13431 6502
rect 13487 6500 13493 6502
rect 13185 6491 13493 6500
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 6089 13032 6190
rect 12990 6080 13046 6089
rect 12990 6015 13046 6024
rect 12636 5506 12756 5534
rect 12176 5234 12204 5506
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 4282 11008 4490
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 9784 3670 9812 4082
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9784 3534 9812 3606
rect 10060 3534 10088 3674
rect 9220 3528 9272 3534
rect 9404 3528 9456 3534
rect 9220 3470 9272 3476
rect 9310 3496 9366 3505
rect 9232 3194 9260 3470
rect 9404 3470 9456 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9310 3431 9366 3440
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8597 2748 8905 2757
rect 8597 2746 8603 2748
rect 8659 2746 8683 2748
rect 8739 2746 8763 2748
rect 8819 2746 8843 2748
rect 8899 2746 8905 2748
rect 8659 2694 8661 2746
rect 8841 2694 8843 2746
rect 8597 2692 8603 2694
rect 8659 2692 8683 2694
rect 8739 2692 8763 2694
rect 8819 2692 8843 2694
rect 8899 2692 8905 2694
rect 8597 2683 8905 2692
rect 8956 2650 8984 2994
rect 9324 2990 9352 3431
rect 9416 3398 9444 3470
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3058 9444 3334
rect 9692 3194 9720 3470
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 10060 2854 10088 3470
rect 10126 3292 10434 3301
rect 10126 3290 10132 3292
rect 10188 3290 10212 3292
rect 10268 3290 10292 3292
rect 10348 3290 10372 3292
rect 10428 3290 10434 3292
rect 10188 3238 10190 3290
rect 10370 3238 10372 3290
rect 10126 3236 10132 3238
rect 10188 3236 10212 3238
rect 10268 3236 10292 3238
rect 10348 3236 10372 3238
rect 10428 3236 10434 3238
rect 10126 3227 10434 3236
rect 10520 2990 10548 3946
rect 10704 3738 10732 4014
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10796 3618 10824 3878
rect 10888 3738 10916 4082
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10796 3590 10916 3618
rect 10888 3534 10916 3590
rect 10980 3534 11008 4218
rect 11072 4214 11100 4422
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11164 3602 11192 4558
rect 11256 4078 11284 5102
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11532 4690 11560 4966
rect 11656 4924 11964 4933
rect 11656 4922 11662 4924
rect 11718 4922 11742 4924
rect 11798 4922 11822 4924
rect 11878 4922 11902 4924
rect 11958 4922 11964 4924
rect 11718 4870 11720 4922
rect 11900 4870 11902 4922
rect 11656 4868 11662 4870
rect 11718 4868 11742 4870
rect 11798 4868 11822 4870
rect 11878 4868 11902 4870
rect 11958 4868 11964 4870
rect 11656 4859 11964 4868
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 12176 4554 12204 4966
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 4282 11376 4422
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11656 3836 11964 3845
rect 11656 3834 11662 3836
rect 11718 3834 11742 3836
rect 11798 3834 11822 3836
rect 11878 3834 11902 3836
rect 11958 3834 11964 3836
rect 11718 3782 11720 3834
rect 11900 3782 11902 3834
rect 11656 3780 11662 3782
rect 11718 3780 11742 3782
rect 11798 3780 11822 3782
rect 11878 3780 11902 3782
rect 11958 3780 11964 3782
rect 11656 3771 11964 3780
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10888 2922 10916 3470
rect 12084 3194 12112 3878
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 3194 12204 3334
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12452 3058 12480 5102
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12544 3194 12572 3470
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 10336 2514 10364 2790
rect 11656 2748 11964 2757
rect 11656 2746 11662 2748
rect 11718 2746 11742 2748
rect 11798 2746 11822 2748
rect 11878 2746 11902 2748
rect 11958 2746 11964 2748
rect 11718 2694 11720 2746
rect 11900 2694 11902 2746
rect 11656 2692 11662 2694
rect 11718 2692 11742 2694
rect 11798 2692 11822 2694
rect 11878 2692 11902 2694
rect 11958 2692 11964 2694
rect 11656 2683 11964 2692
rect 12728 2650 12756 5506
rect 13185 5468 13493 5477
rect 13185 5466 13191 5468
rect 13247 5466 13271 5468
rect 13327 5466 13351 5468
rect 13407 5466 13431 5468
rect 13487 5466 13493 5468
rect 13247 5414 13249 5466
rect 13429 5414 13431 5466
rect 13185 5412 13191 5414
rect 13247 5412 13271 5414
rect 13327 5412 13351 5414
rect 13407 5412 13431 5414
rect 13487 5412 13493 5414
rect 13185 5403 13493 5412
rect 13185 4380 13493 4389
rect 13185 4378 13191 4380
rect 13247 4378 13271 4380
rect 13327 4378 13351 4380
rect 13407 4378 13431 4380
rect 13487 4378 13493 4380
rect 13247 4326 13249 4378
rect 13429 4326 13431 4378
rect 13185 4324 13191 4326
rect 13247 4324 13271 4326
rect 13327 4324 13351 4326
rect 13407 4324 13431 4326
rect 13487 4324 13493 4326
rect 13185 4315 13493 4324
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3738 12940 4082
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13185 3292 13493 3301
rect 13185 3290 13191 3292
rect 13247 3290 13271 3292
rect 13327 3290 13351 3292
rect 13407 3290 13431 3292
rect 13487 3290 13493 3292
rect 13247 3238 13249 3290
rect 13429 3238 13431 3290
rect 13185 3236 13191 3238
rect 13247 3236 13271 3238
rect 13327 3236 13351 3238
rect 13407 3236 13431 3238
rect 13487 3236 13493 3238
rect 13185 3227 13493 3236
rect 13452 3052 13504 3058
rect 13504 3012 13584 3040
rect 13452 2994 13504 3000
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 2596 2440 2648 2446
rect 4160 2440 4212 2446
rect 2596 2382 2648 2388
rect 3896 2388 4160 2394
rect 3896 2382 4212 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 952 800 980 2382
rect 2608 1306 2636 2382
rect 2516 1278 2636 1306
rect 3896 2366 4200 2382
rect 3896 1306 3924 2366
rect 4008 2204 4316 2213
rect 4008 2202 4014 2204
rect 4070 2202 4094 2204
rect 4150 2202 4174 2204
rect 4230 2202 4254 2204
rect 4310 2202 4316 2204
rect 4070 2150 4072 2202
rect 4252 2150 4254 2202
rect 4008 2148 4014 2150
rect 4070 2148 4094 2150
rect 4150 2148 4174 2150
rect 4230 2148 4254 2150
rect 4310 2148 4316 2150
rect 4008 2139 4316 2148
rect 5736 1306 5764 2382
rect 7067 2204 7375 2213
rect 7067 2202 7073 2204
rect 7129 2202 7153 2204
rect 7209 2202 7233 2204
rect 7289 2202 7313 2204
rect 7369 2202 7375 2204
rect 7129 2150 7131 2202
rect 7311 2150 7313 2202
rect 7067 2148 7073 2150
rect 7129 2148 7153 2150
rect 7209 2148 7233 2150
rect 7289 2148 7313 2150
rect 7369 2148 7375 2150
rect 7067 2139 7375 2148
rect 3896 1278 4108 1306
rect 2516 800 2544 1278
rect 4080 800 4108 1278
rect 5644 1278 5764 1306
rect 5644 800 5672 1278
rect 7208 870 7328 898
rect 7208 800 7236 870
rect 938 0 994 800
rect 2502 0 2558 800
rect 4066 0 4122 800
rect 5630 0 5686 800
rect 7194 0 7250 800
rect 7300 762 7328 870
rect 7484 762 7512 2382
rect 8772 800 8800 2382
rect 10126 2204 10434 2213
rect 10126 2202 10132 2204
rect 10188 2202 10212 2204
rect 10268 2202 10292 2204
rect 10348 2202 10372 2204
rect 10428 2202 10434 2204
rect 10188 2150 10190 2202
rect 10370 2150 10372 2202
rect 10126 2148 10132 2150
rect 10188 2148 10212 2150
rect 10268 2148 10292 2150
rect 10348 2148 10372 2150
rect 10428 2148 10434 2150
rect 10126 2139 10434 2148
rect 10336 870 10456 898
rect 10336 800 10364 870
rect 7300 734 7512 762
rect 8758 0 8814 800
rect 10322 0 10378 800
rect 10428 762 10456 870
rect 10612 762 10640 2382
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 11900 800 11928 2314
rect 13004 2009 13032 2314
rect 13185 2204 13493 2213
rect 13185 2202 13191 2204
rect 13247 2202 13271 2204
rect 13327 2202 13351 2204
rect 13407 2202 13431 2204
rect 13487 2202 13493 2204
rect 13247 2150 13249 2202
rect 13429 2150 13431 2202
rect 13185 2148 13191 2150
rect 13247 2148 13271 2150
rect 13327 2148 13351 2150
rect 13407 2148 13431 2150
rect 13487 2148 13493 2150
rect 13185 2139 13493 2148
rect 12990 2000 13046 2009
rect 12990 1935 13046 1944
rect 13556 1578 13584 3012
rect 13464 1550 13584 1578
rect 13464 800 13492 1550
rect 10428 734 10640 762
rect 11886 0 11942 800
rect 13450 0 13506 800
<< via2 >>
rect 4014 14170 4070 14172
rect 4094 14170 4150 14172
rect 4174 14170 4230 14172
rect 4254 14170 4310 14172
rect 4014 14118 4060 14170
rect 4060 14118 4070 14170
rect 4094 14118 4124 14170
rect 4124 14118 4136 14170
rect 4136 14118 4150 14170
rect 4174 14118 4188 14170
rect 4188 14118 4200 14170
rect 4200 14118 4230 14170
rect 4254 14118 4264 14170
rect 4264 14118 4310 14170
rect 4014 14116 4070 14118
rect 4094 14116 4150 14118
rect 4174 14116 4230 14118
rect 4254 14116 4310 14118
rect 7073 14170 7129 14172
rect 7153 14170 7209 14172
rect 7233 14170 7289 14172
rect 7313 14170 7369 14172
rect 7073 14118 7119 14170
rect 7119 14118 7129 14170
rect 7153 14118 7183 14170
rect 7183 14118 7195 14170
rect 7195 14118 7209 14170
rect 7233 14118 7247 14170
rect 7247 14118 7259 14170
rect 7259 14118 7289 14170
rect 7313 14118 7323 14170
rect 7323 14118 7369 14170
rect 7073 14116 7129 14118
rect 7153 14116 7209 14118
rect 7233 14116 7289 14118
rect 7313 14116 7369 14118
rect 10132 14170 10188 14172
rect 10212 14170 10268 14172
rect 10292 14170 10348 14172
rect 10372 14170 10428 14172
rect 10132 14118 10178 14170
rect 10178 14118 10188 14170
rect 10212 14118 10242 14170
rect 10242 14118 10254 14170
rect 10254 14118 10268 14170
rect 10292 14118 10306 14170
rect 10306 14118 10318 14170
rect 10318 14118 10348 14170
rect 10372 14118 10382 14170
rect 10382 14118 10428 14170
rect 10132 14116 10188 14118
rect 10212 14116 10268 14118
rect 10292 14116 10348 14118
rect 10372 14116 10428 14118
rect 13191 14170 13247 14172
rect 13271 14170 13327 14172
rect 13351 14170 13407 14172
rect 13431 14170 13487 14172
rect 13191 14118 13237 14170
rect 13237 14118 13247 14170
rect 13271 14118 13301 14170
rect 13301 14118 13313 14170
rect 13313 14118 13327 14170
rect 13351 14118 13365 14170
rect 13365 14118 13377 14170
rect 13377 14118 13407 14170
rect 13431 14118 13441 14170
rect 13441 14118 13487 14170
rect 13191 14116 13247 14118
rect 13271 14116 13327 14118
rect 13351 14116 13407 14118
rect 13431 14116 13487 14118
rect 13266 13948 13268 13968
rect 13268 13948 13320 13968
rect 13320 13948 13322 13968
rect 13266 13912 13322 13948
rect 2485 13626 2541 13628
rect 2565 13626 2621 13628
rect 2645 13626 2701 13628
rect 2725 13626 2781 13628
rect 2485 13574 2531 13626
rect 2531 13574 2541 13626
rect 2565 13574 2595 13626
rect 2595 13574 2607 13626
rect 2607 13574 2621 13626
rect 2645 13574 2659 13626
rect 2659 13574 2671 13626
rect 2671 13574 2701 13626
rect 2725 13574 2735 13626
rect 2735 13574 2781 13626
rect 2485 13572 2541 13574
rect 2565 13572 2621 13574
rect 2645 13572 2701 13574
rect 2725 13572 2781 13574
rect 5544 13626 5600 13628
rect 5624 13626 5680 13628
rect 5704 13626 5760 13628
rect 5784 13626 5840 13628
rect 5544 13574 5590 13626
rect 5590 13574 5600 13626
rect 5624 13574 5654 13626
rect 5654 13574 5666 13626
rect 5666 13574 5680 13626
rect 5704 13574 5718 13626
rect 5718 13574 5730 13626
rect 5730 13574 5760 13626
rect 5784 13574 5794 13626
rect 5794 13574 5840 13626
rect 5544 13572 5600 13574
rect 5624 13572 5680 13574
rect 5704 13572 5760 13574
rect 5784 13572 5840 13574
rect 4014 13082 4070 13084
rect 4094 13082 4150 13084
rect 4174 13082 4230 13084
rect 4254 13082 4310 13084
rect 4014 13030 4060 13082
rect 4060 13030 4070 13082
rect 4094 13030 4124 13082
rect 4124 13030 4136 13082
rect 4136 13030 4150 13082
rect 4174 13030 4188 13082
rect 4188 13030 4200 13082
rect 4200 13030 4230 13082
rect 4254 13030 4264 13082
rect 4264 13030 4310 13082
rect 4014 13028 4070 13030
rect 4094 13028 4150 13030
rect 4174 13028 4230 13030
rect 4254 13028 4310 13030
rect 2485 12538 2541 12540
rect 2565 12538 2621 12540
rect 2645 12538 2701 12540
rect 2725 12538 2781 12540
rect 2485 12486 2531 12538
rect 2531 12486 2541 12538
rect 2565 12486 2595 12538
rect 2595 12486 2607 12538
rect 2607 12486 2621 12538
rect 2645 12486 2659 12538
rect 2659 12486 2671 12538
rect 2671 12486 2701 12538
rect 2725 12486 2735 12538
rect 2735 12486 2781 12538
rect 2485 12484 2541 12486
rect 2565 12484 2621 12486
rect 2645 12484 2701 12486
rect 2725 12484 2781 12486
rect 4066 12280 4122 12336
rect 4014 11994 4070 11996
rect 4094 11994 4150 11996
rect 4174 11994 4230 11996
rect 4254 11994 4310 11996
rect 4014 11942 4060 11994
rect 4060 11942 4070 11994
rect 4094 11942 4124 11994
rect 4124 11942 4136 11994
rect 4136 11942 4150 11994
rect 4174 11942 4188 11994
rect 4188 11942 4200 11994
rect 4200 11942 4230 11994
rect 4254 11942 4264 11994
rect 4264 11942 4310 11994
rect 4014 11940 4070 11942
rect 4094 11940 4150 11942
rect 4174 11940 4230 11942
rect 4254 11940 4310 11942
rect 2485 11450 2541 11452
rect 2565 11450 2621 11452
rect 2645 11450 2701 11452
rect 2725 11450 2781 11452
rect 2485 11398 2531 11450
rect 2531 11398 2541 11450
rect 2565 11398 2595 11450
rect 2595 11398 2607 11450
rect 2607 11398 2621 11450
rect 2645 11398 2659 11450
rect 2659 11398 2671 11450
rect 2671 11398 2701 11450
rect 2725 11398 2735 11450
rect 2735 11398 2781 11450
rect 2485 11396 2541 11398
rect 2565 11396 2621 11398
rect 2645 11396 2701 11398
rect 2725 11396 2781 11398
rect 4014 10906 4070 10908
rect 4094 10906 4150 10908
rect 4174 10906 4230 10908
rect 4254 10906 4310 10908
rect 4014 10854 4060 10906
rect 4060 10854 4070 10906
rect 4094 10854 4124 10906
rect 4124 10854 4136 10906
rect 4136 10854 4150 10906
rect 4174 10854 4188 10906
rect 4188 10854 4200 10906
rect 4200 10854 4230 10906
rect 4254 10854 4264 10906
rect 4264 10854 4310 10906
rect 4014 10852 4070 10854
rect 4094 10852 4150 10854
rect 4174 10852 4230 10854
rect 4254 10852 4310 10854
rect 2485 10362 2541 10364
rect 2565 10362 2621 10364
rect 2645 10362 2701 10364
rect 2725 10362 2781 10364
rect 2485 10310 2531 10362
rect 2531 10310 2541 10362
rect 2565 10310 2595 10362
rect 2595 10310 2607 10362
rect 2607 10310 2621 10362
rect 2645 10310 2659 10362
rect 2659 10310 2671 10362
rect 2671 10310 2701 10362
rect 2725 10310 2735 10362
rect 2735 10310 2781 10362
rect 2485 10308 2541 10310
rect 2565 10308 2621 10310
rect 2645 10308 2701 10310
rect 2725 10308 2781 10310
rect 5544 12538 5600 12540
rect 5624 12538 5680 12540
rect 5704 12538 5760 12540
rect 5784 12538 5840 12540
rect 5544 12486 5590 12538
rect 5590 12486 5600 12538
rect 5624 12486 5654 12538
rect 5654 12486 5666 12538
rect 5666 12486 5680 12538
rect 5704 12486 5718 12538
rect 5718 12486 5730 12538
rect 5730 12486 5760 12538
rect 5784 12486 5794 12538
rect 5794 12486 5840 12538
rect 5544 12484 5600 12486
rect 5624 12484 5680 12486
rect 5704 12484 5760 12486
rect 5784 12484 5840 12486
rect 5544 11450 5600 11452
rect 5624 11450 5680 11452
rect 5704 11450 5760 11452
rect 5784 11450 5840 11452
rect 5544 11398 5590 11450
rect 5590 11398 5600 11450
rect 5624 11398 5654 11450
rect 5654 11398 5666 11450
rect 5666 11398 5680 11450
rect 5704 11398 5718 11450
rect 5718 11398 5730 11450
rect 5730 11398 5760 11450
rect 5784 11398 5794 11450
rect 5794 11398 5840 11450
rect 5544 11396 5600 11398
rect 5624 11396 5680 11398
rect 5704 11396 5760 11398
rect 5784 11396 5840 11398
rect 2485 9274 2541 9276
rect 2565 9274 2621 9276
rect 2645 9274 2701 9276
rect 2725 9274 2781 9276
rect 2485 9222 2531 9274
rect 2531 9222 2541 9274
rect 2565 9222 2595 9274
rect 2595 9222 2607 9274
rect 2607 9222 2621 9274
rect 2645 9222 2659 9274
rect 2659 9222 2671 9274
rect 2671 9222 2701 9274
rect 2725 9222 2735 9274
rect 2735 9222 2781 9274
rect 2485 9220 2541 9222
rect 2565 9220 2621 9222
rect 2645 9220 2701 9222
rect 2725 9220 2781 9222
rect 4014 9818 4070 9820
rect 4094 9818 4150 9820
rect 4174 9818 4230 9820
rect 4254 9818 4310 9820
rect 4014 9766 4060 9818
rect 4060 9766 4070 9818
rect 4094 9766 4124 9818
rect 4124 9766 4136 9818
rect 4136 9766 4150 9818
rect 4174 9766 4188 9818
rect 4188 9766 4200 9818
rect 4200 9766 4230 9818
rect 4254 9766 4264 9818
rect 4264 9766 4310 9818
rect 4014 9764 4070 9766
rect 4094 9764 4150 9766
rect 4174 9764 4230 9766
rect 4254 9764 4310 9766
rect 5544 10362 5600 10364
rect 5624 10362 5680 10364
rect 5704 10362 5760 10364
rect 5784 10362 5840 10364
rect 5544 10310 5590 10362
rect 5590 10310 5600 10362
rect 5624 10310 5654 10362
rect 5654 10310 5666 10362
rect 5666 10310 5680 10362
rect 5704 10310 5718 10362
rect 5718 10310 5730 10362
rect 5730 10310 5760 10362
rect 5784 10310 5794 10362
rect 5794 10310 5840 10362
rect 5544 10308 5600 10310
rect 5624 10308 5680 10310
rect 5704 10308 5760 10310
rect 5784 10308 5840 10310
rect 938 4120 994 4176
rect 2485 8186 2541 8188
rect 2565 8186 2621 8188
rect 2645 8186 2701 8188
rect 2725 8186 2781 8188
rect 2485 8134 2531 8186
rect 2531 8134 2541 8186
rect 2565 8134 2595 8186
rect 2595 8134 2607 8186
rect 2607 8134 2621 8186
rect 2645 8134 2659 8186
rect 2659 8134 2671 8186
rect 2671 8134 2701 8186
rect 2725 8134 2735 8186
rect 2735 8134 2781 8186
rect 2485 8132 2541 8134
rect 2565 8132 2621 8134
rect 2645 8132 2701 8134
rect 2725 8132 2781 8134
rect 2485 7098 2541 7100
rect 2565 7098 2621 7100
rect 2645 7098 2701 7100
rect 2725 7098 2781 7100
rect 2485 7046 2531 7098
rect 2531 7046 2541 7098
rect 2565 7046 2595 7098
rect 2595 7046 2607 7098
rect 2607 7046 2621 7098
rect 2645 7046 2659 7098
rect 2659 7046 2671 7098
rect 2671 7046 2701 7098
rect 2725 7046 2735 7098
rect 2735 7046 2781 7098
rect 2485 7044 2541 7046
rect 2565 7044 2621 7046
rect 2645 7044 2701 7046
rect 2725 7044 2781 7046
rect 4014 8730 4070 8732
rect 4094 8730 4150 8732
rect 4174 8730 4230 8732
rect 4254 8730 4310 8732
rect 4014 8678 4060 8730
rect 4060 8678 4070 8730
rect 4094 8678 4124 8730
rect 4124 8678 4136 8730
rect 4136 8678 4150 8730
rect 4174 8678 4188 8730
rect 4188 8678 4200 8730
rect 4200 8678 4230 8730
rect 4254 8678 4264 8730
rect 4264 8678 4310 8730
rect 4014 8676 4070 8678
rect 4094 8676 4150 8678
rect 4174 8676 4230 8678
rect 4254 8676 4310 8678
rect 2485 6010 2541 6012
rect 2565 6010 2621 6012
rect 2645 6010 2701 6012
rect 2725 6010 2781 6012
rect 2485 5958 2531 6010
rect 2531 5958 2541 6010
rect 2565 5958 2595 6010
rect 2595 5958 2607 6010
rect 2607 5958 2621 6010
rect 2645 5958 2659 6010
rect 2659 5958 2671 6010
rect 2671 5958 2701 6010
rect 2725 5958 2735 6010
rect 2735 5958 2781 6010
rect 2485 5956 2541 5958
rect 2565 5956 2621 5958
rect 2645 5956 2701 5958
rect 2725 5956 2781 5958
rect 2485 4922 2541 4924
rect 2565 4922 2621 4924
rect 2645 4922 2701 4924
rect 2725 4922 2781 4924
rect 2485 4870 2531 4922
rect 2531 4870 2541 4922
rect 2565 4870 2595 4922
rect 2595 4870 2607 4922
rect 2607 4870 2621 4922
rect 2645 4870 2659 4922
rect 2659 4870 2671 4922
rect 2671 4870 2701 4922
rect 2725 4870 2735 4922
rect 2735 4870 2781 4922
rect 2485 4868 2541 4870
rect 2565 4868 2621 4870
rect 2645 4868 2701 4870
rect 2725 4868 2781 4870
rect 4014 7642 4070 7644
rect 4094 7642 4150 7644
rect 4174 7642 4230 7644
rect 4254 7642 4310 7644
rect 4014 7590 4060 7642
rect 4060 7590 4070 7642
rect 4094 7590 4124 7642
rect 4124 7590 4136 7642
rect 4136 7590 4150 7642
rect 4174 7590 4188 7642
rect 4188 7590 4200 7642
rect 4200 7590 4230 7642
rect 4254 7590 4264 7642
rect 4264 7590 4310 7642
rect 4014 7588 4070 7590
rect 4094 7588 4150 7590
rect 4174 7588 4230 7590
rect 4254 7588 4310 7590
rect 4014 6554 4070 6556
rect 4094 6554 4150 6556
rect 4174 6554 4230 6556
rect 4254 6554 4310 6556
rect 4014 6502 4060 6554
rect 4060 6502 4070 6554
rect 4094 6502 4124 6554
rect 4124 6502 4136 6554
rect 4136 6502 4150 6554
rect 4174 6502 4188 6554
rect 4188 6502 4200 6554
rect 4200 6502 4230 6554
rect 4254 6502 4264 6554
rect 4264 6502 4310 6554
rect 4014 6500 4070 6502
rect 4094 6500 4150 6502
rect 4174 6500 4230 6502
rect 4254 6500 4310 6502
rect 4014 5466 4070 5468
rect 4094 5466 4150 5468
rect 4174 5466 4230 5468
rect 4254 5466 4310 5468
rect 4014 5414 4060 5466
rect 4060 5414 4070 5466
rect 4094 5414 4124 5466
rect 4124 5414 4136 5466
rect 4136 5414 4150 5466
rect 4174 5414 4188 5466
rect 4188 5414 4200 5466
rect 4200 5414 4230 5466
rect 4254 5414 4264 5466
rect 4264 5414 4310 5466
rect 4014 5412 4070 5414
rect 4094 5412 4150 5414
rect 4174 5412 4230 5414
rect 4254 5412 4310 5414
rect 2485 3834 2541 3836
rect 2565 3834 2621 3836
rect 2645 3834 2701 3836
rect 2725 3834 2781 3836
rect 2485 3782 2531 3834
rect 2531 3782 2541 3834
rect 2565 3782 2595 3834
rect 2595 3782 2607 3834
rect 2607 3782 2621 3834
rect 2645 3782 2659 3834
rect 2659 3782 2671 3834
rect 2671 3782 2701 3834
rect 2725 3782 2735 3834
rect 2735 3782 2781 3834
rect 2485 3780 2541 3782
rect 2565 3780 2621 3782
rect 2645 3780 2701 3782
rect 2725 3780 2781 3782
rect 4014 4378 4070 4380
rect 4094 4378 4150 4380
rect 4174 4378 4230 4380
rect 4254 4378 4310 4380
rect 4014 4326 4060 4378
rect 4060 4326 4070 4378
rect 4094 4326 4124 4378
rect 4124 4326 4136 4378
rect 4136 4326 4150 4378
rect 4174 4326 4188 4378
rect 4188 4326 4200 4378
rect 4200 4326 4230 4378
rect 4254 4326 4264 4378
rect 4264 4326 4310 4378
rect 4014 4324 4070 4326
rect 4094 4324 4150 4326
rect 4174 4324 4230 4326
rect 4254 4324 4310 4326
rect 2485 2746 2541 2748
rect 2565 2746 2621 2748
rect 2645 2746 2701 2748
rect 2725 2746 2781 2748
rect 2485 2694 2531 2746
rect 2531 2694 2541 2746
rect 2565 2694 2595 2746
rect 2595 2694 2607 2746
rect 2607 2694 2621 2746
rect 2645 2694 2659 2746
rect 2659 2694 2671 2746
rect 2671 2694 2701 2746
rect 2725 2694 2735 2746
rect 2735 2694 2781 2746
rect 2485 2692 2541 2694
rect 2565 2692 2621 2694
rect 2645 2692 2701 2694
rect 2725 2692 2781 2694
rect 4014 3290 4070 3292
rect 4094 3290 4150 3292
rect 4174 3290 4230 3292
rect 4254 3290 4310 3292
rect 4014 3238 4060 3290
rect 4060 3238 4070 3290
rect 4094 3238 4124 3290
rect 4124 3238 4136 3290
rect 4136 3238 4150 3290
rect 4174 3238 4188 3290
rect 4188 3238 4200 3290
rect 4200 3238 4230 3290
rect 4254 3238 4264 3290
rect 4264 3238 4310 3290
rect 4014 3236 4070 3238
rect 4094 3236 4150 3238
rect 4174 3236 4230 3238
rect 4254 3236 4310 3238
rect 5544 9274 5600 9276
rect 5624 9274 5680 9276
rect 5704 9274 5760 9276
rect 5784 9274 5840 9276
rect 5544 9222 5590 9274
rect 5590 9222 5600 9274
rect 5624 9222 5654 9274
rect 5654 9222 5666 9274
rect 5666 9222 5680 9274
rect 5704 9222 5718 9274
rect 5718 9222 5730 9274
rect 5730 9222 5760 9274
rect 5784 9222 5794 9274
rect 5794 9222 5840 9274
rect 5544 9220 5600 9222
rect 5624 9220 5680 9222
rect 5704 9220 5760 9222
rect 5784 9220 5840 9222
rect 5544 8186 5600 8188
rect 5624 8186 5680 8188
rect 5704 8186 5760 8188
rect 5784 8186 5840 8188
rect 5544 8134 5590 8186
rect 5590 8134 5600 8186
rect 5624 8134 5654 8186
rect 5654 8134 5666 8186
rect 5666 8134 5680 8186
rect 5704 8134 5718 8186
rect 5718 8134 5730 8186
rect 5730 8134 5760 8186
rect 5784 8134 5794 8186
rect 5794 8134 5840 8186
rect 5544 8132 5600 8134
rect 5624 8132 5680 8134
rect 5704 8132 5760 8134
rect 5784 8132 5840 8134
rect 5544 7098 5600 7100
rect 5624 7098 5680 7100
rect 5704 7098 5760 7100
rect 5784 7098 5840 7100
rect 5544 7046 5590 7098
rect 5590 7046 5600 7098
rect 5624 7046 5654 7098
rect 5654 7046 5666 7098
rect 5666 7046 5680 7098
rect 5704 7046 5718 7098
rect 5718 7046 5730 7098
rect 5730 7046 5760 7098
rect 5784 7046 5794 7098
rect 5794 7046 5840 7098
rect 5544 7044 5600 7046
rect 5624 7044 5680 7046
rect 5704 7044 5760 7046
rect 5784 7044 5840 7046
rect 5544 6010 5600 6012
rect 5624 6010 5680 6012
rect 5704 6010 5760 6012
rect 5784 6010 5840 6012
rect 5544 5958 5590 6010
rect 5590 5958 5600 6010
rect 5624 5958 5654 6010
rect 5654 5958 5666 6010
rect 5666 5958 5680 6010
rect 5704 5958 5718 6010
rect 5718 5958 5730 6010
rect 5730 5958 5760 6010
rect 5784 5958 5794 6010
rect 5794 5958 5840 6010
rect 5544 5956 5600 5958
rect 5624 5956 5680 5958
rect 5704 5956 5760 5958
rect 5784 5956 5840 5958
rect 8603 13626 8659 13628
rect 8683 13626 8739 13628
rect 8763 13626 8819 13628
rect 8843 13626 8899 13628
rect 8603 13574 8649 13626
rect 8649 13574 8659 13626
rect 8683 13574 8713 13626
rect 8713 13574 8725 13626
rect 8725 13574 8739 13626
rect 8763 13574 8777 13626
rect 8777 13574 8789 13626
rect 8789 13574 8819 13626
rect 8843 13574 8853 13626
rect 8853 13574 8899 13626
rect 8603 13572 8659 13574
rect 8683 13572 8739 13574
rect 8763 13572 8819 13574
rect 8843 13572 8899 13574
rect 7073 13082 7129 13084
rect 7153 13082 7209 13084
rect 7233 13082 7289 13084
rect 7313 13082 7369 13084
rect 7073 13030 7119 13082
rect 7119 13030 7129 13082
rect 7153 13030 7183 13082
rect 7183 13030 7195 13082
rect 7195 13030 7209 13082
rect 7233 13030 7247 13082
rect 7247 13030 7259 13082
rect 7259 13030 7289 13082
rect 7313 13030 7323 13082
rect 7323 13030 7369 13082
rect 7073 13028 7129 13030
rect 7153 13028 7209 13030
rect 7233 13028 7289 13030
rect 7313 13028 7369 13030
rect 8022 12280 8078 12336
rect 8603 12538 8659 12540
rect 8683 12538 8739 12540
rect 8763 12538 8819 12540
rect 8843 12538 8899 12540
rect 8603 12486 8649 12538
rect 8649 12486 8659 12538
rect 8683 12486 8713 12538
rect 8713 12486 8725 12538
rect 8725 12486 8739 12538
rect 8763 12486 8777 12538
rect 8777 12486 8789 12538
rect 8789 12486 8819 12538
rect 8843 12486 8853 12538
rect 8853 12486 8899 12538
rect 8603 12484 8659 12486
rect 8683 12484 8739 12486
rect 8763 12484 8819 12486
rect 8843 12484 8899 12486
rect 10132 13082 10188 13084
rect 10212 13082 10268 13084
rect 10292 13082 10348 13084
rect 10372 13082 10428 13084
rect 10132 13030 10178 13082
rect 10178 13030 10188 13082
rect 10212 13030 10242 13082
rect 10242 13030 10254 13082
rect 10254 13030 10268 13082
rect 10292 13030 10306 13082
rect 10306 13030 10318 13082
rect 10318 13030 10348 13082
rect 10372 13030 10382 13082
rect 10382 13030 10428 13082
rect 10132 13028 10188 13030
rect 10212 13028 10268 13030
rect 10292 13028 10348 13030
rect 10372 13028 10428 13030
rect 7073 11994 7129 11996
rect 7153 11994 7209 11996
rect 7233 11994 7289 11996
rect 7313 11994 7369 11996
rect 7073 11942 7119 11994
rect 7119 11942 7129 11994
rect 7153 11942 7183 11994
rect 7183 11942 7195 11994
rect 7195 11942 7209 11994
rect 7233 11942 7247 11994
rect 7247 11942 7259 11994
rect 7259 11942 7289 11994
rect 7313 11942 7323 11994
rect 7323 11942 7369 11994
rect 7073 11940 7129 11942
rect 7153 11940 7209 11942
rect 7233 11940 7289 11942
rect 7313 11940 7369 11942
rect 7073 10906 7129 10908
rect 7153 10906 7209 10908
rect 7233 10906 7289 10908
rect 7313 10906 7369 10908
rect 7073 10854 7119 10906
rect 7119 10854 7129 10906
rect 7153 10854 7183 10906
rect 7183 10854 7195 10906
rect 7195 10854 7209 10906
rect 7233 10854 7247 10906
rect 7247 10854 7259 10906
rect 7259 10854 7289 10906
rect 7313 10854 7323 10906
rect 7323 10854 7369 10906
rect 7073 10852 7129 10854
rect 7153 10852 7209 10854
rect 7233 10852 7289 10854
rect 7313 10852 7369 10854
rect 7073 9818 7129 9820
rect 7153 9818 7209 9820
rect 7233 9818 7289 9820
rect 7313 9818 7369 9820
rect 7073 9766 7119 9818
rect 7119 9766 7129 9818
rect 7153 9766 7183 9818
rect 7183 9766 7195 9818
rect 7195 9766 7209 9818
rect 7233 9766 7247 9818
rect 7247 9766 7259 9818
rect 7259 9766 7289 9818
rect 7313 9766 7323 9818
rect 7323 9766 7369 9818
rect 7073 9764 7129 9766
rect 7153 9764 7209 9766
rect 7233 9764 7289 9766
rect 7313 9764 7369 9766
rect 8603 11450 8659 11452
rect 8683 11450 8739 11452
rect 8763 11450 8819 11452
rect 8843 11450 8899 11452
rect 8603 11398 8649 11450
rect 8649 11398 8659 11450
rect 8683 11398 8713 11450
rect 8713 11398 8725 11450
rect 8725 11398 8739 11450
rect 8763 11398 8777 11450
rect 8777 11398 8789 11450
rect 8789 11398 8819 11450
rect 8843 11398 8853 11450
rect 8853 11398 8899 11450
rect 8603 11396 8659 11398
rect 8683 11396 8739 11398
rect 8763 11396 8819 11398
rect 8843 11396 8899 11398
rect 7073 8730 7129 8732
rect 7153 8730 7209 8732
rect 7233 8730 7289 8732
rect 7313 8730 7369 8732
rect 7073 8678 7119 8730
rect 7119 8678 7129 8730
rect 7153 8678 7183 8730
rect 7183 8678 7195 8730
rect 7195 8678 7209 8730
rect 7233 8678 7247 8730
rect 7247 8678 7259 8730
rect 7259 8678 7289 8730
rect 7313 8678 7323 8730
rect 7323 8678 7369 8730
rect 7073 8676 7129 8678
rect 7153 8676 7209 8678
rect 7233 8676 7289 8678
rect 7313 8676 7369 8678
rect 7073 7642 7129 7644
rect 7153 7642 7209 7644
rect 7233 7642 7289 7644
rect 7313 7642 7369 7644
rect 7073 7590 7119 7642
rect 7119 7590 7129 7642
rect 7153 7590 7183 7642
rect 7183 7590 7195 7642
rect 7195 7590 7209 7642
rect 7233 7590 7247 7642
rect 7247 7590 7259 7642
rect 7259 7590 7289 7642
rect 7313 7590 7323 7642
rect 7323 7590 7369 7642
rect 7073 7588 7129 7590
rect 7153 7588 7209 7590
rect 7233 7588 7289 7590
rect 7313 7588 7369 7590
rect 7073 6554 7129 6556
rect 7153 6554 7209 6556
rect 7233 6554 7289 6556
rect 7313 6554 7369 6556
rect 7073 6502 7119 6554
rect 7119 6502 7129 6554
rect 7153 6502 7183 6554
rect 7183 6502 7195 6554
rect 7195 6502 7209 6554
rect 7233 6502 7247 6554
rect 7247 6502 7259 6554
rect 7259 6502 7289 6554
rect 7313 6502 7323 6554
rect 7323 6502 7369 6554
rect 7073 6500 7129 6502
rect 7153 6500 7209 6502
rect 7233 6500 7289 6502
rect 7313 6500 7369 6502
rect 7073 5466 7129 5468
rect 7153 5466 7209 5468
rect 7233 5466 7289 5468
rect 7313 5466 7369 5468
rect 7073 5414 7119 5466
rect 7119 5414 7129 5466
rect 7153 5414 7183 5466
rect 7183 5414 7195 5466
rect 7195 5414 7209 5466
rect 7233 5414 7247 5466
rect 7247 5414 7259 5466
rect 7259 5414 7289 5466
rect 7313 5414 7323 5466
rect 7323 5414 7369 5466
rect 7073 5412 7129 5414
rect 7153 5412 7209 5414
rect 7233 5412 7289 5414
rect 7313 5412 7369 5414
rect 5544 4922 5600 4924
rect 5624 4922 5680 4924
rect 5704 4922 5760 4924
rect 5784 4922 5840 4924
rect 5544 4870 5590 4922
rect 5590 4870 5600 4922
rect 5624 4870 5654 4922
rect 5654 4870 5666 4922
rect 5666 4870 5680 4922
rect 5704 4870 5718 4922
rect 5718 4870 5730 4922
rect 5730 4870 5760 4922
rect 5784 4870 5794 4922
rect 5794 4870 5840 4922
rect 5544 4868 5600 4870
rect 5624 4868 5680 4870
rect 5704 4868 5760 4870
rect 5784 4868 5840 4870
rect 7073 4378 7129 4380
rect 7153 4378 7209 4380
rect 7233 4378 7289 4380
rect 7313 4378 7369 4380
rect 7073 4326 7119 4378
rect 7119 4326 7129 4378
rect 7153 4326 7183 4378
rect 7183 4326 7195 4378
rect 7195 4326 7209 4378
rect 7233 4326 7247 4378
rect 7247 4326 7259 4378
rect 7259 4326 7289 4378
rect 7313 4326 7323 4378
rect 7323 4326 7369 4378
rect 7073 4324 7129 4326
rect 7153 4324 7209 4326
rect 7233 4324 7289 4326
rect 7313 4324 7369 4326
rect 5544 3834 5600 3836
rect 5624 3834 5680 3836
rect 5704 3834 5760 3836
rect 5784 3834 5840 3836
rect 5544 3782 5590 3834
rect 5590 3782 5600 3834
rect 5624 3782 5654 3834
rect 5654 3782 5666 3834
rect 5666 3782 5680 3834
rect 5704 3782 5718 3834
rect 5718 3782 5730 3834
rect 5730 3782 5760 3834
rect 5784 3782 5794 3834
rect 5794 3782 5840 3834
rect 5544 3780 5600 3782
rect 5624 3780 5680 3782
rect 5704 3780 5760 3782
rect 5784 3780 5840 3782
rect 6642 4020 6644 4040
rect 6644 4020 6696 4040
rect 6696 4020 6698 4040
rect 6642 3984 6698 4020
rect 5544 2746 5600 2748
rect 5624 2746 5680 2748
rect 5704 2746 5760 2748
rect 5784 2746 5840 2748
rect 5544 2694 5590 2746
rect 5590 2694 5600 2746
rect 5624 2694 5654 2746
rect 5654 2694 5666 2746
rect 5666 2694 5680 2746
rect 5704 2694 5718 2746
rect 5718 2694 5730 2746
rect 5730 2694 5760 2746
rect 5784 2694 5794 2746
rect 5794 2694 5840 2746
rect 5544 2692 5600 2694
rect 5624 2692 5680 2694
rect 5704 2692 5760 2694
rect 5784 2692 5840 2694
rect 8603 10362 8659 10364
rect 8683 10362 8739 10364
rect 8763 10362 8819 10364
rect 8843 10362 8899 10364
rect 8603 10310 8649 10362
rect 8649 10310 8659 10362
rect 8683 10310 8713 10362
rect 8713 10310 8725 10362
rect 8725 10310 8739 10362
rect 8763 10310 8777 10362
rect 8777 10310 8789 10362
rect 8789 10310 8819 10362
rect 8843 10310 8853 10362
rect 8853 10310 8899 10362
rect 8603 10308 8659 10310
rect 8683 10308 8739 10310
rect 8763 10308 8819 10310
rect 8843 10308 8899 10310
rect 10230 12316 10232 12336
rect 10232 12316 10284 12336
rect 10284 12316 10286 12336
rect 10230 12280 10286 12316
rect 10132 11994 10188 11996
rect 10212 11994 10268 11996
rect 10292 11994 10348 11996
rect 10372 11994 10428 11996
rect 10132 11942 10178 11994
rect 10178 11942 10188 11994
rect 10212 11942 10242 11994
rect 10242 11942 10254 11994
rect 10254 11942 10268 11994
rect 10292 11942 10306 11994
rect 10306 11942 10318 11994
rect 10318 11942 10348 11994
rect 10372 11942 10382 11994
rect 10382 11942 10428 11994
rect 10132 11940 10188 11942
rect 10212 11940 10268 11942
rect 10292 11940 10348 11942
rect 10372 11940 10428 11942
rect 10132 10906 10188 10908
rect 10212 10906 10268 10908
rect 10292 10906 10348 10908
rect 10372 10906 10428 10908
rect 10132 10854 10178 10906
rect 10178 10854 10188 10906
rect 10212 10854 10242 10906
rect 10242 10854 10254 10906
rect 10254 10854 10268 10906
rect 10292 10854 10306 10906
rect 10306 10854 10318 10906
rect 10318 10854 10348 10906
rect 10372 10854 10382 10906
rect 10382 10854 10428 10906
rect 10132 10852 10188 10854
rect 10212 10852 10268 10854
rect 10292 10852 10348 10854
rect 10372 10852 10428 10854
rect 10132 9818 10188 9820
rect 10212 9818 10268 9820
rect 10292 9818 10348 9820
rect 10372 9818 10428 9820
rect 10132 9766 10178 9818
rect 10178 9766 10188 9818
rect 10212 9766 10242 9818
rect 10242 9766 10254 9818
rect 10254 9766 10268 9818
rect 10292 9766 10306 9818
rect 10306 9766 10318 9818
rect 10318 9766 10348 9818
rect 10372 9766 10382 9818
rect 10382 9766 10428 9818
rect 10132 9764 10188 9766
rect 10212 9764 10268 9766
rect 10292 9764 10348 9766
rect 10372 9764 10428 9766
rect 11662 13626 11718 13628
rect 11742 13626 11798 13628
rect 11822 13626 11878 13628
rect 11902 13626 11958 13628
rect 11662 13574 11708 13626
rect 11708 13574 11718 13626
rect 11742 13574 11772 13626
rect 11772 13574 11784 13626
rect 11784 13574 11798 13626
rect 11822 13574 11836 13626
rect 11836 13574 11848 13626
rect 11848 13574 11878 13626
rect 11902 13574 11912 13626
rect 11912 13574 11958 13626
rect 11662 13572 11718 13574
rect 11742 13572 11798 13574
rect 11822 13572 11878 13574
rect 11902 13572 11958 13574
rect 11662 12538 11718 12540
rect 11742 12538 11798 12540
rect 11822 12538 11878 12540
rect 11902 12538 11958 12540
rect 11662 12486 11708 12538
rect 11708 12486 11718 12538
rect 11742 12486 11772 12538
rect 11772 12486 11784 12538
rect 11784 12486 11798 12538
rect 11822 12486 11836 12538
rect 11836 12486 11848 12538
rect 11848 12486 11878 12538
rect 11902 12486 11912 12538
rect 11912 12486 11958 12538
rect 11662 12484 11718 12486
rect 11742 12484 11798 12486
rect 11822 12484 11878 12486
rect 11902 12484 11958 12486
rect 13191 13082 13247 13084
rect 13271 13082 13327 13084
rect 13351 13082 13407 13084
rect 13431 13082 13487 13084
rect 13191 13030 13237 13082
rect 13237 13030 13247 13082
rect 13271 13030 13301 13082
rect 13301 13030 13313 13082
rect 13313 13030 13327 13082
rect 13351 13030 13365 13082
rect 13365 13030 13377 13082
rect 13377 13030 13407 13082
rect 13431 13030 13441 13082
rect 13441 13030 13487 13082
rect 13191 13028 13247 13030
rect 13271 13028 13327 13030
rect 13351 13028 13407 13030
rect 13431 13028 13487 13030
rect 13191 11994 13247 11996
rect 13271 11994 13327 11996
rect 13351 11994 13407 11996
rect 13431 11994 13487 11996
rect 13191 11942 13237 11994
rect 13237 11942 13247 11994
rect 13271 11942 13301 11994
rect 13301 11942 13313 11994
rect 13313 11942 13327 11994
rect 13351 11942 13365 11994
rect 13365 11942 13377 11994
rect 13377 11942 13407 11994
rect 13431 11942 13441 11994
rect 13441 11942 13487 11994
rect 13191 11940 13247 11942
rect 13271 11940 13327 11942
rect 13351 11940 13407 11942
rect 13431 11940 13487 11942
rect 11662 11450 11718 11452
rect 11742 11450 11798 11452
rect 11822 11450 11878 11452
rect 11902 11450 11958 11452
rect 11662 11398 11708 11450
rect 11708 11398 11718 11450
rect 11742 11398 11772 11450
rect 11772 11398 11784 11450
rect 11784 11398 11798 11450
rect 11822 11398 11836 11450
rect 11836 11398 11848 11450
rect 11848 11398 11878 11450
rect 11902 11398 11912 11450
rect 11912 11398 11958 11450
rect 11662 11396 11718 11398
rect 11742 11396 11798 11398
rect 11822 11396 11878 11398
rect 11902 11396 11958 11398
rect 11662 10362 11718 10364
rect 11742 10362 11798 10364
rect 11822 10362 11878 10364
rect 11902 10362 11958 10364
rect 11662 10310 11708 10362
rect 11708 10310 11718 10362
rect 11742 10310 11772 10362
rect 11772 10310 11784 10362
rect 11784 10310 11798 10362
rect 11822 10310 11836 10362
rect 11836 10310 11848 10362
rect 11848 10310 11878 10362
rect 11902 10310 11912 10362
rect 11912 10310 11958 10362
rect 11662 10308 11718 10310
rect 11742 10308 11798 10310
rect 11822 10308 11878 10310
rect 11902 10308 11958 10310
rect 8603 9274 8659 9276
rect 8683 9274 8739 9276
rect 8763 9274 8819 9276
rect 8843 9274 8899 9276
rect 8603 9222 8649 9274
rect 8649 9222 8659 9274
rect 8683 9222 8713 9274
rect 8713 9222 8725 9274
rect 8725 9222 8739 9274
rect 8763 9222 8777 9274
rect 8777 9222 8789 9274
rect 8789 9222 8819 9274
rect 8843 9222 8853 9274
rect 8853 9222 8899 9274
rect 8603 9220 8659 9222
rect 8683 9220 8739 9222
rect 8763 9220 8819 9222
rect 8843 9220 8899 9222
rect 10132 8730 10188 8732
rect 10212 8730 10268 8732
rect 10292 8730 10348 8732
rect 10372 8730 10428 8732
rect 10132 8678 10178 8730
rect 10178 8678 10188 8730
rect 10212 8678 10242 8730
rect 10242 8678 10254 8730
rect 10254 8678 10268 8730
rect 10292 8678 10306 8730
rect 10306 8678 10318 8730
rect 10318 8678 10348 8730
rect 10372 8678 10382 8730
rect 10382 8678 10428 8730
rect 10132 8676 10188 8678
rect 10212 8676 10268 8678
rect 10292 8676 10348 8678
rect 10372 8676 10428 8678
rect 11662 9274 11718 9276
rect 11742 9274 11798 9276
rect 11822 9274 11878 9276
rect 11902 9274 11958 9276
rect 11662 9222 11708 9274
rect 11708 9222 11718 9274
rect 11742 9222 11772 9274
rect 11772 9222 11784 9274
rect 11784 9222 11798 9274
rect 11822 9222 11836 9274
rect 11836 9222 11848 9274
rect 11848 9222 11878 9274
rect 11902 9222 11912 9274
rect 11912 9222 11958 9274
rect 11662 9220 11718 9222
rect 11742 9220 11798 9222
rect 11822 9220 11878 9222
rect 11902 9220 11958 9222
rect 13191 10906 13247 10908
rect 13271 10906 13327 10908
rect 13351 10906 13407 10908
rect 13431 10906 13487 10908
rect 13191 10854 13237 10906
rect 13237 10854 13247 10906
rect 13271 10854 13301 10906
rect 13301 10854 13313 10906
rect 13313 10854 13327 10906
rect 13351 10854 13365 10906
rect 13365 10854 13377 10906
rect 13377 10854 13407 10906
rect 13431 10854 13441 10906
rect 13441 10854 13487 10906
rect 13191 10852 13247 10854
rect 13271 10852 13327 10854
rect 13351 10852 13407 10854
rect 13431 10852 13487 10854
rect 12990 10104 13046 10160
rect 13191 9818 13247 9820
rect 13271 9818 13327 9820
rect 13351 9818 13407 9820
rect 13431 9818 13487 9820
rect 13191 9766 13237 9818
rect 13237 9766 13247 9818
rect 13271 9766 13301 9818
rect 13301 9766 13313 9818
rect 13313 9766 13327 9818
rect 13351 9766 13365 9818
rect 13365 9766 13377 9818
rect 13377 9766 13407 9818
rect 13431 9766 13441 9818
rect 13441 9766 13487 9818
rect 13191 9764 13247 9766
rect 13271 9764 13327 9766
rect 13351 9764 13407 9766
rect 13431 9764 13487 9766
rect 8603 8186 8659 8188
rect 8683 8186 8739 8188
rect 8763 8186 8819 8188
rect 8843 8186 8899 8188
rect 8603 8134 8649 8186
rect 8649 8134 8659 8186
rect 8683 8134 8713 8186
rect 8713 8134 8725 8186
rect 8725 8134 8739 8186
rect 8763 8134 8777 8186
rect 8777 8134 8789 8186
rect 8789 8134 8819 8186
rect 8843 8134 8853 8186
rect 8853 8134 8899 8186
rect 8603 8132 8659 8134
rect 8683 8132 8739 8134
rect 8763 8132 8819 8134
rect 8843 8132 8899 8134
rect 11662 8186 11718 8188
rect 11742 8186 11798 8188
rect 11822 8186 11878 8188
rect 11902 8186 11958 8188
rect 11662 8134 11708 8186
rect 11708 8134 11718 8186
rect 11742 8134 11772 8186
rect 11772 8134 11784 8186
rect 11784 8134 11798 8186
rect 11822 8134 11836 8186
rect 11836 8134 11848 8186
rect 11848 8134 11878 8186
rect 11902 8134 11912 8186
rect 11912 8134 11958 8186
rect 11662 8132 11718 8134
rect 11742 8132 11798 8134
rect 11822 8132 11878 8134
rect 11902 8132 11958 8134
rect 8603 7098 8659 7100
rect 8683 7098 8739 7100
rect 8763 7098 8819 7100
rect 8843 7098 8899 7100
rect 8603 7046 8649 7098
rect 8649 7046 8659 7098
rect 8683 7046 8713 7098
rect 8713 7046 8725 7098
rect 8725 7046 8739 7098
rect 8763 7046 8777 7098
rect 8777 7046 8789 7098
rect 8789 7046 8819 7098
rect 8843 7046 8853 7098
rect 8853 7046 8899 7098
rect 8603 7044 8659 7046
rect 8683 7044 8739 7046
rect 8763 7044 8819 7046
rect 8843 7044 8899 7046
rect 8603 6010 8659 6012
rect 8683 6010 8739 6012
rect 8763 6010 8819 6012
rect 8843 6010 8899 6012
rect 8603 5958 8649 6010
rect 8649 5958 8659 6010
rect 8683 5958 8713 6010
rect 8713 5958 8725 6010
rect 8725 5958 8739 6010
rect 8763 5958 8777 6010
rect 8777 5958 8789 6010
rect 8789 5958 8819 6010
rect 8843 5958 8853 6010
rect 8853 5958 8899 6010
rect 8603 5956 8659 5958
rect 8683 5956 8739 5958
rect 8763 5956 8819 5958
rect 8843 5956 8899 5958
rect 10132 7642 10188 7644
rect 10212 7642 10268 7644
rect 10292 7642 10348 7644
rect 10372 7642 10428 7644
rect 10132 7590 10178 7642
rect 10178 7590 10188 7642
rect 10212 7590 10242 7642
rect 10242 7590 10254 7642
rect 10254 7590 10268 7642
rect 10292 7590 10306 7642
rect 10306 7590 10318 7642
rect 10318 7590 10348 7642
rect 10372 7590 10382 7642
rect 10382 7590 10428 7642
rect 10132 7588 10188 7590
rect 10212 7588 10268 7590
rect 10292 7588 10348 7590
rect 10372 7588 10428 7590
rect 10132 6554 10188 6556
rect 10212 6554 10268 6556
rect 10292 6554 10348 6556
rect 10372 6554 10428 6556
rect 10132 6502 10178 6554
rect 10178 6502 10188 6554
rect 10212 6502 10242 6554
rect 10242 6502 10254 6554
rect 10254 6502 10268 6554
rect 10292 6502 10306 6554
rect 10306 6502 10318 6554
rect 10318 6502 10348 6554
rect 10372 6502 10382 6554
rect 10382 6502 10428 6554
rect 10132 6500 10188 6502
rect 10212 6500 10268 6502
rect 10292 6500 10348 6502
rect 10372 6500 10428 6502
rect 10132 5466 10188 5468
rect 10212 5466 10268 5468
rect 10292 5466 10348 5468
rect 10372 5466 10428 5468
rect 10132 5414 10178 5466
rect 10178 5414 10188 5466
rect 10212 5414 10242 5466
rect 10242 5414 10254 5466
rect 10254 5414 10268 5466
rect 10292 5414 10306 5466
rect 10306 5414 10318 5466
rect 10318 5414 10348 5466
rect 10372 5414 10382 5466
rect 10382 5414 10428 5466
rect 10132 5412 10188 5414
rect 10212 5412 10268 5414
rect 10292 5412 10348 5414
rect 10372 5412 10428 5414
rect 8603 4922 8659 4924
rect 8683 4922 8739 4924
rect 8763 4922 8819 4924
rect 8843 4922 8899 4924
rect 8603 4870 8649 4922
rect 8649 4870 8659 4922
rect 8683 4870 8713 4922
rect 8713 4870 8725 4922
rect 8725 4870 8739 4922
rect 8763 4870 8777 4922
rect 8777 4870 8789 4922
rect 8789 4870 8819 4922
rect 8843 4870 8853 4922
rect 8853 4870 8899 4922
rect 8603 4868 8659 4870
rect 8683 4868 8739 4870
rect 8763 4868 8819 4870
rect 8843 4868 8899 4870
rect 11662 7098 11718 7100
rect 11742 7098 11798 7100
rect 11822 7098 11878 7100
rect 11902 7098 11958 7100
rect 11662 7046 11708 7098
rect 11708 7046 11718 7098
rect 11742 7046 11772 7098
rect 11772 7046 11784 7098
rect 11784 7046 11798 7098
rect 11822 7046 11836 7098
rect 11836 7046 11848 7098
rect 11848 7046 11878 7098
rect 11902 7046 11912 7098
rect 11912 7046 11958 7098
rect 11662 7044 11718 7046
rect 11742 7044 11798 7046
rect 11822 7044 11878 7046
rect 11902 7044 11958 7046
rect 7194 3576 7250 3632
rect 7010 3440 7066 3496
rect 7838 3440 7894 3496
rect 7073 3290 7129 3292
rect 7153 3290 7209 3292
rect 7233 3290 7289 3292
rect 7313 3290 7369 3292
rect 7073 3238 7119 3290
rect 7119 3238 7129 3290
rect 7153 3238 7183 3290
rect 7183 3238 7195 3290
rect 7195 3238 7209 3290
rect 7233 3238 7247 3290
rect 7247 3238 7259 3290
rect 7259 3238 7289 3290
rect 7313 3238 7323 3290
rect 7323 3238 7369 3290
rect 7073 3236 7129 3238
rect 7153 3236 7209 3238
rect 7233 3236 7289 3238
rect 7313 3236 7369 3238
rect 9126 3984 9182 4040
rect 8603 3834 8659 3836
rect 8683 3834 8739 3836
rect 8763 3834 8819 3836
rect 8843 3834 8899 3836
rect 8603 3782 8649 3834
rect 8649 3782 8659 3834
rect 8683 3782 8713 3834
rect 8713 3782 8725 3834
rect 8725 3782 8739 3834
rect 8763 3782 8777 3834
rect 8777 3782 8789 3834
rect 8789 3782 8819 3834
rect 8843 3782 8853 3834
rect 8853 3782 8899 3834
rect 8603 3780 8659 3782
rect 8683 3780 8739 3782
rect 8763 3780 8819 3782
rect 8843 3780 8899 3782
rect 8390 3576 8446 3632
rect 9034 3596 9090 3632
rect 9034 3576 9036 3596
rect 9036 3576 9088 3596
rect 9088 3576 9090 3596
rect 8482 3440 8538 3496
rect 10132 4378 10188 4380
rect 10212 4378 10268 4380
rect 10292 4378 10348 4380
rect 10372 4378 10428 4380
rect 10132 4326 10178 4378
rect 10178 4326 10188 4378
rect 10212 4326 10242 4378
rect 10242 4326 10254 4378
rect 10254 4326 10268 4378
rect 10292 4326 10306 4378
rect 10306 4326 10318 4378
rect 10318 4326 10348 4378
rect 10372 4326 10382 4378
rect 10382 4326 10428 4378
rect 10132 4324 10188 4326
rect 10212 4324 10268 4326
rect 10292 4324 10348 4326
rect 10372 4324 10428 4326
rect 11662 6010 11718 6012
rect 11742 6010 11798 6012
rect 11822 6010 11878 6012
rect 11902 6010 11958 6012
rect 11662 5958 11708 6010
rect 11708 5958 11718 6010
rect 11742 5958 11772 6010
rect 11772 5958 11784 6010
rect 11784 5958 11798 6010
rect 11822 5958 11836 6010
rect 11836 5958 11848 6010
rect 11848 5958 11878 6010
rect 11902 5958 11912 6010
rect 11912 5958 11958 6010
rect 11662 5956 11718 5958
rect 11742 5956 11798 5958
rect 11822 5956 11878 5958
rect 11902 5956 11958 5958
rect 13191 8730 13247 8732
rect 13271 8730 13327 8732
rect 13351 8730 13407 8732
rect 13431 8730 13487 8732
rect 13191 8678 13237 8730
rect 13237 8678 13247 8730
rect 13271 8678 13301 8730
rect 13301 8678 13313 8730
rect 13313 8678 13327 8730
rect 13351 8678 13365 8730
rect 13365 8678 13377 8730
rect 13377 8678 13407 8730
rect 13431 8678 13441 8730
rect 13441 8678 13487 8730
rect 13191 8676 13247 8678
rect 13271 8676 13327 8678
rect 13351 8676 13407 8678
rect 13431 8676 13487 8678
rect 13191 7642 13247 7644
rect 13271 7642 13327 7644
rect 13351 7642 13407 7644
rect 13431 7642 13487 7644
rect 13191 7590 13237 7642
rect 13237 7590 13247 7642
rect 13271 7590 13301 7642
rect 13301 7590 13313 7642
rect 13313 7590 13327 7642
rect 13351 7590 13365 7642
rect 13365 7590 13377 7642
rect 13377 7590 13407 7642
rect 13431 7590 13441 7642
rect 13441 7590 13487 7642
rect 13191 7588 13247 7590
rect 13271 7588 13327 7590
rect 13351 7588 13407 7590
rect 13431 7588 13487 7590
rect 13191 6554 13247 6556
rect 13271 6554 13327 6556
rect 13351 6554 13407 6556
rect 13431 6554 13487 6556
rect 13191 6502 13237 6554
rect 13237 6502 13247 6554
rect 13271 6502 13301 6554
rect 13301 6502 13313 6554
rect 13313 6502 13327 6554
rect 13351 6502 13365 6554
rect 13365 6502 13377 6554
rect 13377 6502 13407 6554
rect 13431 6502 13441 6554
rect 13441 6502 13487 6554
rect 13191 6500 13247 6502
rect 13271 6500 13327 6502
rect 13351 6500 13407 6502
rect 13431 6500 13487 6502
rect 12990 6024 13046 6080
rect 9310 3440 9366 3496
rect 8603 2746 8659 2748
rect 8683 2746 8739 2748
rect 8763 2746 8819 2748
rect 8843 2746 8899 2748
rect 8603 2694 8649 2746
rect 8649 2694 8659 2746
rect 8683 2694 8713 2746
rect 8713 2694 8725 2746
rect 8725 2694 8739 2746
rect 8763 2694 8777 2746
rect 8777 2694 8789 2746
rect 8789 2694 8819 2746
rect 8843 2694 8853 2746
rect 8853 2694 8899 2746
rect 8603 2692 8659 2694
rect 8683 2692 8739 2694
rect 8763 2692 8819 2694
rect 8843 2692 8899 2694
rect 10132 3290 10188 3292
rect 10212 3290 10268 3292
rect 10292 3290 10348 3292
rect 10372 3290 10428 3292
rect 10132 3238 10178 3290
rect 10178 3238 10188 3290
rect 10212 3238 10242 3290
rect 10242 3238 10254 3290
rect 10254 3238 10268 3290
rect 10292 3238 10306 3290
rect 10306 3238 10318 3290
rect 10318 3238 10348 3290
rect 10372 3238 10382 3290
rect 10382 3238 10428 3290
rect 10132 3236 10188 3238
rect 10212 3236 10268 3238
rect 10292 3236 10348 3238
rect 10372 3236 10428 3238
rect 11662 4922 11718 4924
rect 11742 4922 11798 4924
rect 11822 4922 11878 4924
rect 11902 4922 11958 4924
rect 11662 4870 11708 4922
rect 11708 4870 11718 4922
rect 11742 4870 11772 4922
rect 11772 4870 11784 4922
rect 11784 4870 11798 4922
rect 11822 4870 11836 4922
rect 11836 4870 11848 4922
rect 11848 4870 11878 4922
rect 11902 4870 11912 4922
rect 11912 4870 11958 4922
rect 11662 4868 11718 4870
rect 11742 4868 11798 4870
rect 11822 4868 11878 4870
rect 11902 4868 11958 4870
rect 11662 3834 11718 3836
rect 11742 3834 11798 3836
rect 11822 3834 11878 3836
rect 11902 3834 11958 3836
rect 11662 3782 11708 3834
rect 11708 3782 11718 3834
rect 11742 3782 11772 3834
rect 11772 3782 11784 3834
rect 11784 3782 11798 3834
rect 11822 3782 11836 3834
rect 11836 3782 11848 3834
rect 11848 3782 11878 3834
rect 11902 3782 11912 3834
rect 11912 3782 11958 3834
rect 11662 3780 11718 3782
rect 11742 3780 11798 3782
rect 11822 3780 11878 3782
rect 11902 3780 11958 3782
rect 11662 2746 11718 2748
rect 11742 2746 11798 2748
rect 11822 2746 11878 2748
rect 11902 2746 11958 2748
rect 11662 2694 11708 2746
rect 11708 2694 11718 2746
rect 11742 2694 11772 2746
rect 11772 2694 11784 2746
rect 11784 2694 11798 2746
rect 11822 2694 11836 2746
rect 11836 2694 11848 2746
rect 11848 2694 11878 2746
rect 11902 2694 11912 2746
rect 11912 2694 11958 2746
rect 11662 2692 11718 2694
rect 11742 2692 11798 2694
rect 11822 2692 11878 2694
rect 11902 2692 11958 2694
rect 13191 5466 13247 5468
rect 13271 5466 13327 5468
rect 13351 5466 13407 5468
rect 13431 5466 13487 5468
rect 13191 5414 13237 5466
rect 13237 5414 13247 5466
rect 13271 5414 13301 5466
rect 13301 5414 13313 5466
rect 13313 5414 13327 5466
rect 13351 5414 13365 5466
rect 13365 5414 13377 5466
rect 13377 5414 13407 5466
rect 13431 5414 13441 5466
rect 13441 5414 13487 5466
rect 13191 5412 13247 5414
rect 13271 5412 13327 5414
rect 13351 5412 13407 5414
rect 13431 5412 13487 5414
rect 13191 4378 13247 4380
rect 13271 4378 13327 4380
rect 13351 4378 13407 4380
rect 13431 4378 13487 4380
rect 13191 4326 13237 4378
rect 13237 4326 13247 4378
rect 13271 4326 13301 4378
rect 13301 4326 13313 4378
rect 13313 4326 13327 4378
rect 13351 4326 13365 4378
rect 13365 4326 13377 4378
rect 13377 4326 13407 4378
rect 13431 4326 13441 4378
rect 13441 4326 13487 4378
rect 13191 4324 13247 4326
rect 13271 4324 13327 4326
rect 13351 4324 13407 4326
rect 13431 4324 13487 4326
rect 13191 3290 13247 3292
rect 13271 3290 13327 3292
rect 13351 3290 13407 3292
rect 13431 3290 13487 3292
rect 13191 3238 13237 3290
rect 13237 3238 13247 3290
rect 13271 3238 13301 3290
rect 13301 3238 13313 3290
rect 13313 3238 13327 3290
rect 13351 3238 13365 3290
rect 13365 3238 13377 3290
rect 13377 3238 13407 3290
rect 13431 3238 13441 3290
rect 13441 3238 13487 3290
rect 13191 3236 13247 3238
rect 13271 3236 13327 3238
rect 13351 3236 13407 3238
rect 13431 3236 13487 3238
rect 4014 2202 4070 2204
rect 4094 2202 4150 2204
rect 4174 2202 4230 2204
rect 4254 2202 4310 2204
rect 4014 2150 4060 2202
rect 4060 2150 4070 2202
rect 4094 2150 4124 2202
rect 4124 2150 4136 2202
rect 4136 2150 4150 2202
rect 4174 2150 4188 2202
rect 4188 2150 4200 2202
rect 4200 2150 4230 2202
rect 4254 2150 4264 2202
rect 4264 2150 4310 2202
rect 4014 2148 4070 2150
rect 4094 2148 4150 2150
rect 4174 2148 4230 2150
rect 4254 2148 4310 2150
rect 7073 2202 7129 2204
rect 7153 2202 7209 2204
rect 7233 2202 7289 2204
rect 7313 2202 7369 2204
rect 7073 2150 7119 2202
rect 7119 2150 7129 2202
rect 7153 2150 7183 2202
rect 7183 2150 7195 2202
rect 7195 2150 7209 2202
rect 7233 2150 7247 2202
rect 7247 2150 7259 2202
rect 7259 2150 7289 2202
rect 7313 2150 7323 2202
rect 7323 2150 7369 2202
rect 7073 2148 7129 2150
rect 7153 2148 7209 2150
rect 7233 2148 7289 2150
rect 7313 2148 7369 2150
rect 10132 2202 10188 2204
rect 10212 2202 10268 2204
rect 10292 2202 10348 2204
rect 10372 2202 10428 2204
rect 10132 2150 10178 2202
rect 10178 2150 10188 2202
rect 10212 2150 10242 2202
rect 10242 2150 10254 2202
rect 10254 2150 10268 2202
rect 10292 2150 10306 2202
rect 10306 2150 10318 2202
rect 10318 2150 10348 2202
rect 10372 2150 10382 2202
rect 10382 2150 10428 2202
rect 10132 2148 10188 2150
rect 10212 2148 10268 2150
rect 10292 2148 10348 2150
rect 10372 2148 10428 2150
rect 13191 2202 13247 2204
rect 13271 2202 13327 2204
rect 13351 2202 13407 2204
rect 13431 2202 13487 2204
rect 13191 2150 13237 2202
rect 13237 2150 13247 2202
rect 13271 2150 13301 2202
rect 13301 2150 13313 2202
rect 13313 2150 13327 2202
rect 13351 2150 13365 2202
rect 13365 2150 13377 2202
rect 13377 2150 13407 2202
rect 13431 2150 13441 2202
rect 13441 2150 13487 2202
rect 13191 2148 13247 2150
rect 13271 2148 13327 2150
rect 13351 2148 13407 2150
rect 13431 2148 13487 2150
rect 12990 1944 13046 2000
<< metal3 >>
rect 4004 14176 4320 14177
rect 4004 14112 4010 14176
rect 4074 14112 4090 14176
rect 4154 14112 4170 14176
rect 4234 14112 4250 14176
rect 4314 14112 4320 14176
rect 4004 14111 4320 14112
rect 7063 14176 7379 14177
rect 7063 14112 7069 14176
rect 7133 14112 7149 14176
rect 7213 14112 7229 14176
rect 7293 14112 7309 14176
rect 7373 14112 7379 14176
rect 7063 14111 7379 14112
rect 10122 14176 10438 14177
rect 10122 14112 10128 14176
rect 10192 14112 10208 14176
rect 10272 14112 10288 14176
rect 10352 14112 10368 14176
rect 10432 14112 10438 14176
rect 10122 14111 10438 14112
rect 13181 14176 13497 14177
rect 13181 14112 13187 14176
rect 13251 14112 13267 14176
rect 13331 14112 13347 14176
rect 13411 14112 13427 14176
rect 13491 14112 13497 14176
rect 13657 14152 14457 14272
rect 13181 14111 13497 14112
rect 13261 13970 13327 13973
rect 13678 13970 13738 14152
rect 13261 13968 13738 13970
rect 13261 13912 13266 13968
rect 13322 13912 13738 13968
rect 13261 13910 13738 13912
rect 13261 13907 13327 13910
rect 2475 13632 2791 13633
rect 2475 13568 2481 13632
rect 2545 13568 2561 13632
rect 2625 13568 2641 13632
rect 2705 13568 2721 13632
rect 2785 13568 2791 13632
rect 2475 13567 2791 13568
rect 5534 13632 5850 13633
rect 5534 13568 5540 13632
rect 5604 13568 5620 13632
rect 5684 13568 5700 13632
rect 5764 13568 5780 13632
rect 5844 13568 5850 13632
rect 5534 13567 5850 13568
rect 8593 13632 8909 13633
rect 8593 13568 8599 13632
rect 8663 13568 8679 13632
rect 8743 13568 8759 13632
rect 8823 13568 8839 13632
rect 8903 13568 8909 13632
rect 8593 13567 8909 13568
rect 11652 13632 11968 13633
rect 11652 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11898 13632
rect 11962 13568 11968 13632
rect 11652 13567 11968 13568
rect 4004 13088 4320 13089
rect 4004 13024 4010 13088
rect 4074 13024 4090 13088
rect 4154 13024 4170 13088
rect 4234 13024 4250 13088
rect 4314 13024 4320 13088
rect 4004 13023 4320 13024
rect 7063 13088 7379 13089
rect 7063 13024 7069 13088
rect 7133 13024 7149 13088
rect 7213 13024 7229 13088
rect 7293 13024 7309 13088
rect 7373 13024 7379 13088
rect 7063 13023 7379 13024
rect 10122 13088 10438 13089
rect 10122 13024 10128 13088
rect 10192 13024 10208 13088
rect 10272 13024 10288 13088
rect 10352 13024 10368 13088
rect 10432 13024 10438 13088
rect 10122 13023 10438 13024
rect 13181 13088 13497 13089
rect 13181 13024 13187 13088
rect 13251 13024 13267 13088
rect 13331 13024 13347 13088
rect 13411 13024 13427 13088
rect 13491 13024 13497 13088
rect 13181 13023 13497 13024
rect 2475 12544 2791 12545
rect 2475 12480 2481 12544
rect 2545 12480 2561 12544
rect 2625 12480 2641 12544
rect 2705 12480 2721 12544
rect 2785 12480 2791 12544
rect 2475 12479 2791 12480
rect 5534 12544 5850 12545
rect 5534 12480 5540 12544
rect 5604 12480 5620 12544
rect 5684 12480 5700 12544
rect 5764 12480 5780 12544
rect 5844 12480 5850 12544
rect 5534 12479 5850 12480
rect 8593 12544 8909 12545
rect 8593 12480 8599 12544
rect 8663 12480 8679 12544
rect 8743 12480 8759 12544
rect 8823 12480 8839 12544
rect 8903 12480 8909 12544
rect 8593 12479 8909 12480
rect 11652 12544 11968 12545
rect 11652 12480 11658 12544
rect 11722 12480 11738 12544
rect 11802 12480 11818 12544
rect 11882 12480 11898 12544
rect 11962 12480 11968 12544
rect 11652 12479 11968 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 8017 12338 8083 12341
rect 10225 12338 10291 12341
rect 8017 12336 10291 12338
rect 8017 12280 8022 12336
rect 8078 12280 10230 12336
rect 10286 12280 10291 12336
rect 8017 12278 10291 12280
rect 8017 12275 8083 12278
rect 10225 12275 10291 12278
rect 4004 12000 4320 12001
rect 4004 11936 4010 12000
rect 4074 11936 4090 12000
rect 4154 11936 4170 12000
rect 4234 11936 4250 12000
rect 4314 11936 4320 12000
rect 4004 11935 4320 11936
rect 7063 12000 7379 12001
rect 7063 11936 7069 12000
rect 7133 11936 7149 12000
rect 7213 11936 7229 12000
rect 7293 11936 7309 12000
rect 7373 11936 7379 12000
rect 7063 11935 7379 11936
rect 10122 12000 10438 12001
rect 10122 11936 10128 12000
rect 10192 11936 10208 12000
rect 10272 11936 10288 12000
rect 10352 11936 10368 12000
rect 10432 11936 10438 12000
rect 10122 11935 10438 11936
rect 13181 12000 13497 12001
rect 13181 11936 13187 12000
rect 13251 11936 13267 12000
rect 13331 11936 13347 12000
rect 13411 11936 13427 12000
rect 13491 11936 13497 12000
rect 13181 11935 13497 11936
rect 2475 11456 2791 11457
rect 2475 11392 2481 11456
rect 2545 11392 2561 11456
rect 2625 11392 2641 11456
rect 2705 11392 2721 11456
rect 2785 11392 2791 11456
rect 2475 11391 2791 11392
rect 5534 11456 5850 11457
rect 5534 11392 5540 11456
rect 5604 11392 5620 11456
rect 5684 11392 5700 11456
rect 5764 11392 5780 11456
rect 5844 11392 5850 11456
rect 5534 11391 5850 11392
rect 8593 11456 8909 11457
rect 8593 11392 8599 11456
rect 8663 11392 8679 11456
rect 8743 11392 8759 11456
rect 8823 11392 8839 11456
rect 8903 11392 8909 11456
rect 8593 11391 8909 11392
rect 11652 11456 11968 11457
rect 11652 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11898 11456
rect 11962 11392 11968 11456
rect 11652 11391 11968 11392
rect 4004 10912 4320 10913
rect 4004 10848 4010 10912
rect 4074 10848 4090 10912
rect 4154 10848 4170 10912
rect 4234 10848 4250 10912
rect 4314 10848 4320 10912
rect 4004 10847 4320 10848
rect 7063 10912 7379 10913
rect 7063 10848 7069 10912
rect 7133 10848 7149 10912
rect 7213 10848 7229 10912
rect 7293 10848 7309 10912
rect 7373 10848 7379 10912
rect 7063 10847 7379 10848
rect 10122 10912 10438 10913
rect 10122 10848 10128 10912
rect 10192 10848 10208 10912
rect 10272 10848 10288 10912
rect 10352 10848 10368 10912
rect 10432 10848 10438 10912
rect 10122 10847 10438 10848
rect 13181 10912 13497 10913
rect 13181 10848 13187 10912
rect 13251 10848 13267 10912
rect 13331 10848 13347 10912
rect 13411 10848 13427 10912
rect 13491 10848 13497 10912
rect 13181 10847 13497 10848
rect 2475 10368 2791 10369
rect 2475 10304 2481 10368
rect 2545 10304 2561 10368
rect 2625 10304 2641 10368
rect 2705 10304 2721 10368
rect 2785 10304 2791 10368
rect 2475 10303 2791 10304
rect 5534 10368 5850 10369
rect 5534 10304 5540 10368
rect 5604 10304 5620 10368
rect 5684 10304 5700 10368
rect 5764 10304 5780 10368
rect 5844 10304 5850 10368
rect 5534 10303 5850 10304
rect 8593 10368 8909 10369
rect 8593 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8909 10368
rect 8593 10303 8909 10304
rect 11652 10368 11968 10369
rect 11652 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11898 10368
rect 11962 10304 11968 10368
rect 11652 10303 11968 10304
rect 12985 10162 13051 10165
rect 13657 10162 14457 10192
rect 12985 10160 14457 10162
rect 12985 10104 12990 10160
rect 13046 10104 14457 10160
rect 12985 10102 14457 10104
rect 12985 10099 13051 10102
rect 13657 10072 14457 10102
rect 4004 9824 4320 9825
rect 4004 9760 4010 9824
rect 4074 9760 4090 9824
rect 4154 9760 4170 9824
rect 4234 9760 4250 9824
rect 4314 9760 4320 9824
rect 4004 9759 4320 9760
rect 7063 9824 7379 9825
rect 7063 9760 7069 9824
rect 7133 9760 7149 9824
rect 7213 9760 7229 9824
rect 7293 9760 7309 9824
rect 7373 9760 7379 9824
rect 7063 9759 7379 9760
rect 10122 9824 10438 9825
rect 10122 9760 10128 9824
rect 10192 9760 10208 9824
rect 10272 9760 10288 9824
rect 10352 9760 10368 9824
rect 10432 9760 10438 9824
rect 10122 9759 10438 9760
rect 13181 9824 13497 9825
rect 13181 9760 13187 9824
rect 13251 9760 13267 9824
rect 13331 9760 13347 9824
rect 13411 9760 13427 9824
rect 13491 9760 13497 9824
rect 13181 9759 13497 9760
rect 2475 9280 2791 9281
rect 2475 9216 2481 9280
rect 2545 9216 2561 9280
rect 2625 9216 2641 9280
rect 2705 9216 2721 9280
rect 2785 9216 2791 9280
rect 2475 9215 2791 9216
rect 5534 9280 5850 9281
rect 5534 9216 5540 9280
rect 5604 9216 5620 9280
rect 5684 9216 5700 9280
rect 5764 9216 5780 9280
rect 5844 9216 5850 9280
rect 5534 9215 5850 9216
rect 8593 9280 8909 9281
rect 8593 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8909 9280
rect 8593 9215 8909 9216
rect 11652 9280 11968 9281
rect 11652 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11898 9280
rect 11962 9216 11968 9280
rect 11652 9215 11968 9216
rect 4004 8736 4320 8737
rect 4004 8672 4010 8736
rect 4074 8672 4090 8736
rect 4154 8672 4170 8736
rect 4234 8672 4250 8736
rect 4314 8672 4320 8736
rect 4004 8671 4320 8672
rect 7063 8736 7379 8737
rect 7063 8672 7069 8736
rect 7133 8672 7149 8736
rect 7213 8672 7229 8736
rect 7293 8672 7309 8736
rect 7373 8672 7379 8736
rect 7063 8671 7379 8672
rect 10122 8736 10438 8737
rect 10122 8672 10128 8736
rect 10192 8672 10208 8736
rect 10272 8672 10288 8736
rect 10352 8672 10368 8736
rect 10432 8672 10438 8736
rect 10122 8671 10438 8672
rect 13181 8736 13497 8737
rect 13181 8672 13187 8736
rect 13251 8672 13267 8736
rect 13331 8672 13347 8736
rect 13411 8672 13427 8736
rect 13491 8672 13497 8736
rect 13181 8671 13497 8672
rect 2475 8192 2791 8193
rect 2475 8128 2481 8192
rect 2545 8128 2561 8192
rect 2625 8128 2641 8192
rect 2705 8128 2721 8192
rect 2785 8128 2791 8192
rect 2475 8127 2791 8128
rect 5534 8192 5850 8193
rect 5534 8128 5540 8192
rect 5604 8128 5620 8192
rect 5684 8128 5700 8192
rect 5764 8128 5780 8192
rect 5844 8128 5850 8192
rect 5534 8127 5850 8128
rect 8593 8192 8909 8193
rect 8593 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8909 8192
rect 8593 8127 8909 8128
rect 11652 8192 11968 8193
rect 11652 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11898 8192
rect 11962 8128 11968 8192
rect 11652 8127 11968 8128
rect 4004 7648 4320 7649
rect 4004 7584 4010 7648
rect 4074 7584 4090 7648
rect 4154 7584 4170 7648
rect 4234 7584 4250 7648
rect 4314 7584 4320 7648
rect 4004 7583 4320 7584
rect 7063 7648 7379 7649
rect 7063 7584 7069 7648
rect 7133 7584 7149 7648
rect 7213 7584 7229 7648
rect 7293 7584 7309 7648
rect 7373 7584 7379 7648
rect 7063 7583 7379 7584
rect 10122 7648 10438 7649
rect 10122 7584 10128 7648
rect 10192 7584 10208 7648
rect 10272 7584 10288 7648
rect 10352 7584 10368 7648
rect 10432 7584 10438 7648
rect 10122 7583 10438 7584
rect 13181 7648 13497 7649
rect 13181 7584 13187 7648
rect 13251 7584 13267 7648
rect 13331 7584 13347 7648
rect 13411 7584 13427 7648
rect 13491 7584 13497 7648
rect 13181 7583 13497 7584
rect 2475 7104 2791 7105
rect 2475 7040 2481 7104
rect 2545 7040 2561 7104
rect 2625 7040 2641 7104
rect 2705 7040 2721 7104
rect 2785 7040 2791 7104
rect 2475 7039 2791 7040
rect 5534 7104 5850 7105
rect 5534 7040 5540 7104
rect 5604 7040 5620 7104
rect 5684 7040 5700 7104
rect 5764 7040 5780 7104
rect 5844 7040 5850 7104
rect 5534 7039 5850 7040
rect 8593 7104 8909 7105
rect 8593 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8909 7104
rect 8593 7039 8909 7040
rect 11652 7104 11968 7105
rect 11652 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11898 7104
rect 11962 7040 11968 7104
rect 11652 7039 11968 7040
rect 4004 6560 4320 6561
rect 4004 6496 4010 6560
rect 4074 6496 4090 6560
rect 4154 6496 4170 6560
rect 4234 6496 4250 6560
rect 4314 6496 4320 6560
rect 4004 6495 4320 6496
rect 7063 6560 7379 6561
rect 7063 6496 7069 6560
rect 7133 6496 7149 6560
rect 7213 6496 7229 6560
rect 7293 6496 7309 6560
rect 7373 6496 7379 6560
rect 7063 6495 7379 6496
rect 10122 6560 10438 6561
rect 10122 6496 10128 6560
rect 10192 6496 10208 6560
rect 10272 6496 10288 6560
rect 10352 6496 10368 6560
rect 10432 6496 10438 6560
rect 10122 6495 10438 6496
rect 13181 6560 13497 6561
rect 13181 6496 13187 6560
rect 13251 6496 13267 6560
rect 13331 6496 13347 6560
rect 13411 6496 13427 6560
rect 13491 6496 13497 6560
rect 13181 6495 13497 6496
rect 12985 6082 13051 6085
rect 13657 6082 14457 6112
rect 12985 6080 14457 6082
rect 12985 6024 12990 6080
rect 13046 6024 14457 6080
rect 12985 6022 14457 6024
rect 12985 6019 13051 6022
rect 2475 6016 2791 6017
rect 2475 5952 2481 6016
rect 2545 5952 2561 6016
rect 2625 5952 2641 6016
rect 2705 5952 2721 6016
rect 2785 5952 2791 6016
rect 2475 5951 2791 5952
rect 5534 6016 5850 6017
rect 5534 5952 5540 6016
rect 5604 5952 5620 6016
rect 5684 5952 5700 6016
rect 5764 5952 5780 6016
rect 5844 5952 5850 6016
rect 5534 5951 5850 5952
rect 8593 6016 8909 6017
rect 8593 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8909 6016
rect 8593 5951 8909 5952
rect 11652 6016 11968 6017
rect 11652 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11898 6016
rect 11962 5952 11968 6016
rect 13657 5992 14457 6022
rect 11652 5951 11968 5952
rect 4004 5472 4320 5473
rect 4004 5408 4010 5472
rect 4074 5408 4090 5472
rect 4154 5408 4170 5472
rect 4234 5408 4250 5472
rect 4314 5408 4320 5472
rect 4004 5407 4320 5408
rect 7063 5472 7379 5473
rect 7063 5408 7069 5472
rect 7133 5408 7149 5472
rect 7213 5408 7229 5472
rect 7293 5408 7309 5472
rect 7373 5408 7379 5472
rect 7063 5407 7379 5408
rect 10122 5472 10438 5473
rect 10122 5408 10128 5472
rect 10192 5408 10208 5472
rect 10272 5408 10288 5472
rect 10352 5408 10368 5472
rect 10432 5408 10438 5472
rect 10122 5407 10438 5408
rect 13181 5472 13497 5473
rect 13181 5408 13187 5472
rect 13251 5408 13267 5472
rect 13331 5408 13347 5472
rect 13411 5408 13427 5472
rect 13491 5408 13497 5472
rect 13181 5407 13497 5408
rect 2475 4928 2791 4929
rect 2475 4864 2481 4928
rect 2545 4864 2561 4928
rect 2625 4864 2641 4928
rect 2705 4864 2721 4928
rect 2785 4864 2791 4928
rect 2475 4863 2791 4864
rect 5534 4928 5850 4929
rect 5534 4864 5540 4928
rect 5604 4864 5620 4928
rect 5684 4864 5700 4928
rect 5764 4864 5780 4928
rect 5844 4864 5850 4928
rect 5534 4863 5850 4864
rect 8593 4928 8909 4929
rect 8593 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8909 4928
rect 8593 4863 8909 4864
rect 11652 4928 11968 4929
rect 11652 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11898 4928
rect 11962 4864 11968 4928
rect 11652 4863 11968 4864
rect 4004 4384 4320 4385
rect 4004 4320 4010 4384
rect 4074 4320 4090 4384
rect 4154 4320 4170 4384
rect 4234 4320 4250 4384
rect 4314 4320 4320 4384
rect 4004 4319 4320 4320
rect 7063 4384 7379 4385
rect 7063 4320 7069 4384
rect 7133 4320 7149 4384
rect 7213 4320 7229 4384
rect 7293 4320 7309 4384
rect 7373 4320 7379 4384
rect 7063 4319 7379 4320
rect 10122 4384 10438 4385
rect 10122 4320 10128 4384
rect 10192 4320 10208 4384
rect 10272 4320 10288 4384
rect 10352 4320 10368 4384
rect 10432 4320 10438 4384
rect 10122 4319 10438 4320
rect 13181 4384 13497 4385
rect 13181 4320 13187 4384
rect 13251 4320 13267 4384
rect 13331 4320 13347 4384
rect 13411 4320 13427 4384
rect 13491 4320 13497 4384
rect 13181 4319 13497 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 6637 4042 6703 4045
rect 9121 4042 9187 4045
rect 6637 4040 9187 4042
rect 6637 3984 6642 4040
rect 6698 3984 9126 4040
rect 9182 3984 9187 4040
rect 6637 3982 9187 3984
rect 6637 3979 6703 3982
rect 9121 3979 9187 3982
rect 2475 3840 2791 3841
rect 2475 3776 2481 3840
rect 2545 3776 2561 3840
rect 2625 3776 2641 3840
rect 2705 3776 2721 3840
rect 2785 3776 2791 3840
rect 2475 3775 2791 3776
rect 5534 3840 5850 3841
rect 5534 3776 5540 3840
rect 5604 3776 5620 3840
rect 5684 3776 5700 3840
rect 5764 3776 5780 3840
rect 5844 3776 5850 3840
rect 5534 3775 5850 3776
rect 8593 3840 8909 3841
rect 8593 3776 8599 3840
rect 8663 3776 8679 3840
rect 8743 3776 8759 3840
rect 8823 3776 8839 3840
rect 8903 3776 8909 3840
rect 8593 3775 8909 3776
rect 11652 3840 11968 3841
rect 11652 3776 11658 3840
rect 11722 3776 11738 3840
rect 11802 3776 11818 3840
rect 11882 3776 11898 3840
rect 11962 3776 11968 3840
rect 11652 3775 11968 3776
rect 7189 3634 7255 3637
rect 8385 3634 8451 3637
rect 9029 3634 9095 3637
rect 7189 3632 9095 3634
rect 7189 3576 7194 3632
rect 7250 3576 8390 3632
rect 8446 3576 9034 3632
rect 9090 3576 9095 3632
rect 7189 3574 9095 3576
rect 7189 3571 7255 3574
rect 8385 3571 8451 3574
rect 9029 3571 9095 3574
rect 7005 3498 7071 3501
rect 7833 3498 7899 3501
rect 8477 3498 8543 3501
rect 9305 3498 9371 3501
rect 7005 3496 9371 3498
rect 7005 3440 7010 3496
rect 7066 3440 7838 3496
rect 7894 3440 8482 3496
rect 8538 3440 9310 3496
rect 9366 3440 9371 3496
rect 7005 3438 9371 3440
rect 7005 3435 7071 3438
rect 7833 3435 7899 3438
rect 8477 3435 8543 3438
rect 9305 3435 9371 3438
rect 4004 3296 4320 3297
rect 4004 3232 4010 3296
rect 4074 3232 4090 3296
rect 4154 3232 4170 3296
rect 4234 3232 4250 3296
rect 4314 3232 4320 3296
rect 4004 3231 4320 3232
rect 7063 3296 7379 3297
rect 7063 3232 7069 3296
rect 7133 3232 7149 3296
rect 7213 3232 7229 3296
rect 7293 3232 7309 3296
rect 7373 3232 7379 3296
rect 7063 3231 7379 3232
rect 10122 3296 10438 3297
rect 10122 3232 10128 3296
rect 10192 3232 10208 3296
rect 10272 3232 10288 3296
rect 10352 3232 10368 3296
rect 10432 3232 10438 3296
rect 10122 3231 10438 3232
rect 13181 3296 13497 3297
rect 13181 3232 13187 3296
rect 13251 3232 13267 3296
rect 13331 3232 13347 3296
rect 13411 3232 13427 3296
rect 13491 3232 13497 3296
rect 13181 3231 13497 3232
rect 2475 2752 2791 2753
rect 2475 2688 2481 2752
rect 2545 2688 2561 2752
rect 2625 2688 2641 2752
rect 2705 2688 2721 2752
rect 2785 2688 2791 2752
rect 2475 2687 2791 2688
rect 5534 2752 5850 2753
rect 5534 2688 5540 2752
rect 5604 2688 5620 2752
rect 5684 2688 5700 2752
rect 5764 2688 5780 2752
rect 5844 2688 5850 2752
rect 5534 2687 5850 2688
rect 8593 2752 8909 2753
rect 8593 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8909 2752
rect 8593 2687 8909 2688
rect 11652 2752 11968 2753
rect 11652 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11898 2752
rect 11962 2688 11968 2752
rect 11652 2687 11968 2688
rect 4004 2208 4320 2209
rect 4004 2144 4010 2208
rect 4074 2144 4090 2208
rect 4154 2144 4170 2208
rect 4234 2144 4250 2208
rect 4314 2144 4320 2208
rect 4004 2143 4320 2144
rect 7063 2208 7379 2209
rect 7063 2144 7069 2208
rect 7133 2144 7149 2208
rect 7213 2144 7229 2208
rect 7293 2144 7309 2208
rect 7373 2144 7379 2208
rect 7063 2143 7379 2144
rect 10122 2208 10438 2209
rect 10122 2144 10128 2208
rect 10192 2144 10208 2208
rect 10272 2144 10288 2208
rect 10352 2144 10368 2208
rect 10432 2144 10438 2208
rect 10122 2143 10438 2144
rect 13181 2208 13497 2209
rect 13181 2144 13187 2208
rect 13251 2144 13267 2208
rect 13331 2144 13347 2208
rect 13411 2144 13427 2208
rect 13491 2144 13497 2208
rect 13181 2143 13497 2144
rect 12985 2002 13051 2005
rect 13657 2002 14457 2032
rect 12985 2000 14457 2002
rect 12985 1944 12990 2000
rect 13046 1944 14457 2000
rect 12985 1942 14457 1944
rect 12985 1939 13051 1942
rect 13657 1912 14457 1942
<< via3 >>
rect 4010 14172 4074 14176
rect 4010 14116 4014 14172
rect 4014 14116 4070 14172
rect 4070 14116 4074 14172
rect 4010 14112 4074 14116
rect 4090 14172 4154 14176
rect 4090 14116 4094 14172
rect 4094 14116 4150 14172
rect 4150 14116 4154 14172
rect 4090 14112 4154 14116
rect 4170 14172 4234 14176
rect 4170 14116 4174 14172
rect 4174 14116 4230 14172
rect 4230 14116 4234 14172
rect 4170 14112 4234 14116
rect 4250 14172 4314 14176
rect 4250 14116 4254 14172
rect 4254 14116 4310 14172
rect 4310 14116 4314 14172
rect 4250 14112 4314 14116
rect 7069 14172 7133 14176
rect 7069 14116 7073 14172
rect 7073 14116 7129 14172
rect 7129 14116 7133 14172
rect 7069 14112 7133 14116
rect 7149 14172 7213 14176
rect 7149 14116 7153 14172
rect 7153 14116 7209 14172
rect 7209 14116 7213 14172
rect 7149 14112 7213 14116
rect 7229 14172 7293 14176
rect 7229 14116 7233 14172
rect 7233 14116 7289 14172
rect 7289 14116 7293 14172
rect 7229 14112 7293 14116
rect 7309 14172 7373 14176
rect 7309 14116 7313 14172
rect 7313 14116 7369 14172
rect 7369 14116 7373 14172
rect 7309 14112 7373 14116
rect 10128 14172 10192 14176
rect 10128 14116 10132 14172
rect 10132 14116 10188 14172
rect 10188 14116 10192 14172
rect 10128 14112 10192 14116
rect 10208 14172 10272 14176
rect 10208 14116 10212 14172
rect 10212 14116 10268 14172
rect 10268 14116 10272 14172
rect 10208 14112 10272 14116
rect 10288 14172 10352 14176
rect 10288 14116 10292 14172
rect 10292 14116 10348 14172
rect 10348 14116 10352 14172
rect 10288 14112 10352 14116
rect 10368 14172 10432 14176
rect 10368 14116 10372 14172
rect 10372 14116 10428 14172
rect 10428 14116 10432 14172
rect 10368 14112 10432 14116
rect 13187 14172 13251 14176
rect 13187 14116 13191 14172
rect 13191 14116 13247 14172
rect 13247 14116 13251 14172
rect 13187 14112 13251 14116
rect 13267 14172 13331 14176
rect 13267 14116 13271 14172
rect 13271 14116 13327 14172
rect 13327 14116 13331 14172
rect 13267 14112 13331 14116
rect 13347 14172 13411 14176
rect 13347 14116 13351 14172
rect 13351 14116 13407 14172
rect 13407 14116 13411 14172
rect 13347 14112 13411 14116
rect 13427 14172 13491 14176
rect 13427 14116 13431 14172
rect 13431 14116 13487 14172
rect 13487 14116 13491 14172
rect 13427 14112 13491 14116
rect 2481 13628 2545 13632
rect 2481 13572 2485 13628
rect 2485 13572 2541 13628
rect 2541 13572 2545 13628
rect 2481 13568 2545 13572
rect 2561 13628 2625 13632
rect 2561 13572 2565 13628
rect 2565 13572 2621 13628
rect 2621 13572 2625 13628
rect 2561 13568 2625 13572
rect 2641 13628 2705 13632
rect 2641 13572 2645 13628
rect 2645 13572 2701 13628
rect 2701 13572 2705 13628
rect 2641 13568 2705 13572
rect 2721 13628 2785 13632
rect 2721 13572 2725 13628
rect 2725 13572 2781 13628
rect 2781 13572 2785 13628
rect 2721 13568 2785 13572
rect 5540 13628 5604 13632
rect 5540 13572 5544 13628
rect 5544 13572 5600 13628
rect 5600 13572 5604 13628
rect 5540 13568 5604 13572
rect 5620 13628 5684 13632
rect 5620 13572 5624 13628
rect 5624 13572 5680 13628
rect 5680 13572 5684 13628
rect 5620 13568 5684 13572
rect 5700 13628 5764 13632
rect 5700 13572 5704 13628
rect 5704 13572 5760 13628
rect 5760 13572 5764 13628
rect 5700 13568 5764 13572
rect 5780 13628 5844 13632
rect 5780 13572 5784 13628
rect 5784 13572 5840 13628
rect 5840 13572 5844 13628
rect 5780 13568 5844 13572
rect 8599 13628 8663 13632
rect 8599 13572 8603 13628
rect 8603 13572 8659 13628
rect 8659 13572 8663 13628
rect 8599 13568 8663 13572
rect 8679 13628 8743 13632
rect 8679 13572 8683 13628
rect 8683 13572 8739 13628
rect 8739 13572 8743 13628
rect 8679 13568 8743 13572
rect 8759 13628 8823 13632
rect 8759 13572 8763 13628
rect 8763 13572 8819 13628
rect 8819 13572 8823 13628
rect 8759 13568 8823 13572
rect 8839 13628 8903 13632
rect 8839 13572 8843 13628
rect 8843 13572 8899 13628
rect 8899 13572 8903 13628
rect 8839 13568 8903 13572
rect 11658 13628 11722 13632
rect 11658 13572 11662 13628
rect 11662 13572 11718 13628
rect 11718 13572 11722 13628
rect 11658 13568 11722 13572
rect 11738 13628 11802 13632
rect 11738 13572 11742 13628
rect 11742 13572 11798 13628
rect 11798 13572 11802 13628
rect 11738 13568 11802 13572
rect 11818 13628 11882 13632
rect 11818 13572 11822 13628
rect 11822 13572 11878 13628
rect 11878 13572 11882 13628
rect 11818 13568 11882 13572
rect 11898 13628 11962 13632
rect 11898 13572 11902 13628
rect 11902 13572 11958 13628
rect 11958 13572 11962 13628
rect 11898 13568 11962 13572
rect 4010 13084 4074 13088
rect 4010 13028 4014 13084
rect 4014 13028 4070 13084
rect 4070 13028 4074 13084
rect 4010 13024 4074 13028
rect 4090 13084 4154 13088
rect 4090 13028 4094 13084
rect 4094 13028 4150 13084
rect 4150 13028 4154 13084
rect 4090 13024 4154 13028
rect 4170 13084 4234 13088
rect 4170 13028 4174 13084
rect 4174 13028 4230 13084
rect 4230 13028 4234 13084
rect 4170 13024 4234 13028
rect 4250 13084 4314 13088
rect 4250 13028 4254 13084
rect 4254 13028 4310 13084
rect 4310 13028 4314 13084
rect 4250 13024 4314 13028
rect 7069 13084 7133 13088
rect 7069 13028 7073 13084
rect 7073 13028 7129 13084
rect 7129 13028 7133 13084
rect 7069 13024 7133 13028
rect 7149 13084 7213 13088
rect 7149 13028 7153 13084
rect 7153 13028 7209 13084
rect 7209 13028 7213 13084
rect 7149 13024 7213 13028
rect 7229 13084 7293 13088
rect 7229 13028 7233 13084
rect 7233 13028 7289 13084
rect 7289 13028 7293 13084
rect 7229 13024 7293 13028
rect 7309 13084 7373 13088
rect 7309 13028 7313 13084
rect 7313 13028 7369 13084
rect 7369 13028 7373 13084
rect 7309 13024 7373 13028
rect 10128 13084 10192 13088
rect 10128 13028 10132 13084
rect 10132 13028 10188 13084
rect 10188 13028 10192 13084
rect 10128 13024 10192 13028
rect 10208 13084 10272 13088
rect 10208 13028 10212 13084
rect 10212 13028 10268 13084
rect 10268 13028 10272 13084
rect 10208 13024 10272 13028
rect 10288 13084 10352 13088
rect 10288 13028 10292 13084
rect 10292 13028 10348 13084
rect 10348 13028 10352 13084
rect 10288 13024 10352 13028
rect 10368 13084 10432 13088
rect 10368 13028 10372 13084
rect 10372 13028 10428 13084
rect 10428 13028 10432 13084
rect 10368 13024 10432 13028
rect 13187 13084 13251 13088
rect 13187 13028 13191 13084
rect 13191 13028 13247 13084
rect 13247 13028 13251 13084
rect 13187 13024 13251 13028
rect 13267 13084 13331 13088
rect 13267 13028 13271 13084
rect 13271 13028 13327 13084
rect 13327 13028 13331 13084
rect 13267 13024 13331 13028
rect 13347 13084 13411 13088
rect 13347 13028 13351 13084
rect 13351 13028 13407 13084
rect 13407 13028 13411 13084
rect 13347 13024 13411 13028
rect 13427 13084 13491 13088
rect 13427 13028 13431 13084
rect 13431 13028 13487 13084
rect 13487 13028 13491 13084
rect 13427 13024 13491 13028
rect 2481 12540 2545 12544
rect 2481 12484 2485 12540
rect 2485 12484 2541 12540
rect 2541 12484 2545 12540
rect 2481 12480 2545 12484
rect 2561 12540 2625 12544
rect 2561 12484 2565 12540
rect 2565 12484 2621 12540
rect 2621 12484 2625 12540
rect 2561 12480 2625 12484
rect 2641 12540 2705 12544
rect 2641 12484 2645 12540
rect 2645 12484 2701 12540
rect 2701 12484 2705 12540
rect 2641 12480 2705 12484
rect 2721 12540 2785 12544
rect 2721 12484 2725 12540
rect 2725 12484 2781 12540
rect 2781 12484 2785 12540
rect 2721 12480 2785 12484
rect 5540 12540 5604 12544
rect 5540 12484 5544 12540
rect 5544 12484 5600 12540
rect 5600 12484 5604 12540
rect 5540 12480 5604 12484
rect 5620 12540 5684 12544
rect 5620 12484 5624 12540
rect 5624 12484 5680 12540
rect 5680 12484 5684 12540
rect 5620 12480 5684 12484
rect 5700 12540 5764 12544
rect 5700 12484 5704 12540
rect 5704 12484 5760 12540
rect 5760 12484 5764 12540
rect 5700 12480 5764 12484
rect 5780 12540 5844 12544
rect 5780 12484 5784 12540
rect 5784 12484 5840 12540
rect 5840 12484 5844 12540
rect 5780 12480 5844 12484
rect 8599 12540 8663 12544
rect 8599 12484 8603 12540
rect 8603 12484 8659 12540
rect 8659 12484 8663 12540
rect 8599 12480 8663 12484
rect 8679 12540 8743 12544
rect 8679 12484 8683 12540
rect 8683 12484 8739 12540
rect 8739 12484 8743 12540
rect 8679 12480 8743 12484
rect 8759 12540 8823 12544
rect 8759 12484 8763 12540
rect 8763 12484 8819 12540
rect 8819 12484 8823 12540
rect 8759 12480 8823 12484
rect 8839 12540 8903 12544
rect 8839 12484 8843 12540
rect 8843 12484 8899 12540
rect 8899 12484 8903 12540
rect 8839 12480 8903 12484
rect 11658 12540 11722 12544
rect 11658 12484 11662 12540
rect 11662 12484 11718 12540
rect 11718 12484 11722 12540
rect 11658 12480 11722 12484
rect 11738 12540 11802 12544
rect 11738 12484 11742 12540
rect 11742 12484 11798 12540
rect 11798 12484 11802 12540
rect 11738 12480 11802 12484
rect 11818 12540 11882 12544
rect 11818 12484 11822 12540
rect 11822 12484 11878 12540
rect 11878 12484 11882 12540
rect 11818 12480 11882 12484
rect 11898 12540 11962 12544
rect 11898 12484 11902 12540
rect 11902 12484 11958 12540
rect 11958 12484 11962 12540
rect 11898 12480 11962 12484
rect 4010 11996 4074 12000
rect 4010 11940 4014 11996
rect 4014 11940 4070 11996
rect 4070 11940 4074 11996
rect 4010 11936 4074 11940
rect 4090 11996 4154 12000
rect 4090 11940 4094 11996
rect 4094 11940 4150 11996
rect 4150 11940 4154 11996
rect 4090 11936 4154 11940
rect 4170 11996 4234 12000
rect 4170 11940 4174 11996
rect 4174 11940 4230 11996
rect 4230 11940 4234 11996
rect 4170 11936 4234 11940
rect 4250 11996 4314 12000
rect 4250 11940 4254 11996
rect 4254 11940 4310 11996
rect 4310 11940 4314 11996
rect 4250 11936 4314 11940
rect 7069 11996 7133 12000
rect 7069 11940 7073 11996
rect 7073 11940 7129 11996
rect 7129 11940 7133 11996
rect 7069 11936 7133 11940
rect 7149 11996 7213 12000
rect 7149 11940 7153 11996
rect 7153 11940 7209 11996
rect 7209 11940 7213 11996
rect 7149 11936 7213 11940
rect 7229 11996 7293 12000
rect 7229 11940 7233 11996
rect 7233 11940 7289 11996
rect 7289 11940 7293 11996
rect 7229 11936 7293 11940
rect 7309 11996 7373 12000
rect 7309 11940 7313 11996
rect 7313 11940 7369 11996
rect 7369 11940 7373 11996
rect 7309 11936 7373 11940
rect 10128 11996 10192 12000
rect 10128 11940 10132 11996
rect 10132 11940 10188 11996
rect 10188 11940 10192 11996
rect 10128 11936 10192 11940
rect 10208 11996 10272 12000
rect 10208 11940 10212 11996
rect 10212 11940 10268 11996
rect 10268 11940 10272 11996
rect 10208 11936 10272 11940
rect 10288 11996 10352 12000
rect 10288 11940 10292 11996
rect 10292 11940 10348 11996
rect 10348 11940 10352 11996
rect 10288 11936 10352 11940
rect 10368 11996 10432 12000
rect 10368 11940 10372 11996
rect 10372 11940 10428 11996
rect 10428 11940 10432 11996
rect 10368 11936 10432 11940
rect 13187 11996 13251 12000
rect 13187 11940 13191 11996
rect 13191 11940 13247 11996
rect 13247 11940 13251 11996
rect 13187 11936 13251 11940
rect 13267 11996 13331 12000
rect 13267 11940 13271 11996
rect 13271 11940 13327 11996
rect 13327 11940 13331 11996
rect 13267 11936 13331 11940
rect 13347 11996 13411 12000
rect 13347 11940 13351 11996
rect 13351 11940 13407 11996
rect 13407 11940 13411 11996
rect 13347 11936 13411 11940
rect 13427 11996 13491 12000
rect 13427 11940 13431 11996
rect 13431 11940 13487 11996
rect 13487 11940 13491 11996
rect 13427 11936 13491 11940
rect 2481 11452 2545 11456
rect 2481 11396 2485 11452
rect 2485 11396 2541 11452
rect 2541 11396 2545 11452
rect 2481 11392 2545 11396
rect 2561 11452 2625 11456
rect 2561 11396 2565 11452
rect 2565 11396 2621 11452
rect 2621 11396 2625 11452
rect 2561 11392 2625 11396
rect 2641 11452 2705 11456
rect 2641 11396 2645 11452
rect 2645 11396 2701 11452
rect 2701 11396 2705 11452
rect 2641 11392 2705 11396
rect 2721 11452 2785 11456
rect 2721 11396 2725 11452
rect 2725 11396 2781 11452
rect 2781 11396 2785 11452
rect 2721 11392 2785 11396
rect 5540 11452 5604 11456
rect 5540 11396 5544 11452
rect 5544 11396 5600 11452
rect 5600 11396 5604 11452
rect 5540 11392 5604 11396
rect 5620 11452 5684 11456
rect 5620 11396 5624 11452
rect 5624 11396 5680 11452
rect 5680 11396 5684 11452
rect 5620 11392 5684 11396
rect 5700 11452 5764 11456
rect 5700 11396 5704 11452
rect 5704 11396 5760 11452
rect 5760 11396 5764 11452
rect 5700 11392 5764 11396
rect 5780 11452 5844 11456
rect 5780 11396 5784 11452
rect 5784 11396 5840 11452
rect 5840 11396 5844 11452
rect 5780 11392 5844 11396
rect 8599 11452 8663 11456
rect 8599 11396 8603 11452
rect 8603 11396 8659 11452
rect 8659 11396 8663 11452
rect 8599 11392 8663 11396
rect 8679 11452 8743 11456
rect 8679 11396 8683 11452
rect 8683 11396 8739 11452
rect 8739 11396 8743 11452
rect 8679 11392 8743 11396
rect 8759 11452 8823 11456
rect 8759 11396 8763 11452
rect 8763 11396 8819 11452
rect 8819 11396 8823 11452
rect 8759 11392 8823 11396
rect 8839 11452 8903 11456
rect 8839 11396 8843 11452
rect 8843 11396 8899 11452
rect 8899 11396 8903 11452
rect 8839 11392 8903 11396
rect 11658 11452 11722 11456
rect 11658 11396 11662 11452
rect 11662 11396 11718 11452
rect 11718 11396 11722 11452
rect 11658 11392 11722 11396
rect 11738 11452 11802 11456
rect 11738 11396 11742 11452
rect 11742 11396 11798 11452
rect 11798 11396 11802 11452
rect 11738 11392 11802 11396
rect 11818 11452 11882 11456
rect 11818 11396 11822 11452
rect 11822 11396 11878 11452
rect 11878 11396 11882 11452
rect 11818 11392 11882 11396
rect 11898 11452 11962 11456
rect 11898 11396 11902 11452
rect 11902 11396 11958 11452
rect 11958 11396 11962 11452
rect 11898 11392 11962 11396
rect 4010 10908 4074 10912
rect 4010 10852 4014 10908
rect 4014 10852 4070 10908
rect 4070 10852 4074 10908
rect 4010 10848 4074 10852
rect 4090 10908 4154 10912
rect 4090 10852 4094 10908
rect 4094 10852 4150 10908
rect 4150 10852 4154 10908
rect 4090 10848 4154 10852
rect 4170 10908 4234 10912
rect 4170 10852 4174 10908
rect 4174 10852 4230 10908
rect 4230 10852 4234 10908
rect 4170 10848 4234 10852
rect 4250 10908 4314 10912
rect 4250 10852 4254 10908
rect 4254 10852 4310 10908
rect 4310 10852 4314 10908
rect 4250 10848 4314 10852
rect 7069 10908 7133 10912
rect 7069 10852 7073 10908
rect 7073 10852 7129 10908
rect 7129 10852 7133 10908
rect 7069 10848 7133 10852
rect 7149 10908 7213 10912
rect 7149 10852 7153 10908
rect 7153 10852 7209 10908
rect 7209 10852 7213 10908
rect 7149 10848 7213 10852
rect 7229 10908 7293 10912
rect 7229 10852 7233 10908
rect 7233 10852 7289 10908
rect 7289 10852 7293 10908
rect 7229 10848 7293 10852
rect 7309 10908 7373 10912
rect 7309 10852 7313 10908
rect 7313 10852 7369 10908
rect 7369 10852 7373 10908
rect 7309 10848 7373 10852
rect 10128 10908 10192 10912
rect 10128 10852 10132 10908
rect 10132 10852 10188 10908
rect 10188 10852 10192 10908
rect 10128 10848 10192 10852
rect 10208 10908 10272 10912
rect 10208 10852 10212 10908
rect 10212 10852 10268 10908
rect 10268 10852 10272 10908
rect 10208 10848 10272 10852
rect 10288 10908 10352 10912
rect 10288 10852 10292 10908
rect 10292 10852 10348 10908
rect 10348 10852 10352 10908
rect 10288 10848 10352 10852
rect 10368 10908 10432 10912
rect 10368 10852 10372 10908
rect 10372 10852 10428 10908
rect 10428 10852 10432 10908
rect 10368 10848 10432 10852
rect 13187 10908 13251 10912
rect 13187 10852 13191 10908
rect 13191 10852 13247 10908
rect 13247 10852 13251 10908
rect 13187 10848 13251 10852
rect 13267 10908 13331 10912
rect 13267 10852 13271 10908
rect 13271 10852 13327 10908
rect 13327 10852 13331 10908
rect 13267 10848 13331 10852
rect 13347 10908 13411 10912
rect 13347 10852 13351 10908
rect 13351 10852 13407 10908
rect 13407 10852 13411 10908
rect 13347 10848 13411 10852
rect 13427 10908 13491 10912
rect 13427 10852 13431 10908
rect 13431 10852 13487 10908
rect 13487 10852 13491 10908
rect 13427 10848 13491 10852
rect 2481 10364 2545 10368
rect 2481 10308 2485 10364
rect 2485 10308 2541 10364
rect 2541 10308 2545 10364
rect 2481 10304 2545 10308
rect 2561 10364 2625 10368
rect 2561 10308 2565 10364
rect 2565 10308 2621 10364
rect 2621 10308 2625 10364
rect 2561 10304 2625 10308
rect 2641 10364 2705 10368
rect 2641 10308 2645 10364
rect 2645 10308 2701 10364
rect 2701 10308 2705 10364
rect 2641 10304 2705 10308
rect 2721 10364 2785 10368
rect 2721 10308 2725 10364
rect 2725 10308 2781 10364
rect 2781 10308 2785 10364
rect 2721 10304 2785 10308
rect 5540 10364 5604 10368
rect 5540 10308 5544 10364
rect 5544 10308 5600 10364
rect 5600 10308 5604 10364
rect 5540 10304 5604 10308
rect 5620 10364 5684 10368
rect 5620 10308 5624 10364
rect 5624 10308 5680 10364
rect 5680 10308 5684 10364
rect 5620 10304 5684 10308
rect 5700 10364 5764 10368
rect 5700 10308 5704 10364
rect 5704 10308 5760 10364
rect 5760 10308 5764 10364
rect 5700 10304 5764 10308
rect 5780 10364 5844 10368
rect 5780 10308 5784 10364
rect 5784 10308 5840 10364
rect 5840 10308 5844 10364
rect 5780 10304 5844 10308
rect 8599 10364 8663 10368
rect 8599 10308 8603 10364
rect 8603 10308 8659 10364
rect 8659 10308 8663 10364
rect 8599 10304 8663 10308
rect 8679 10364 8743 10368
rect 8679 10308 8683 10364
rect 8683 10308 8739 10364
rect 8739 10308 8743 10364
rect 8679 10304 8743 10308
rect 8759 10364 8823 10368
rect 8759 10308 8763 10364
rect 8763 10308 8819 10364
rect 8819 10308 8823 10364
rect 8759 10304 8823 10308
rect 8839 10364 8903 10368
rect 8839 10308 8843 10364
rect 8843 10308 8899 10364
rect 8899 10308 8903 10364
rect 8839 10304 8903 10308
rect 11658 10364 11722 10368
rect 11658 10308 11662 10364
rect 11662 10308 11718 10364
rect 11718 10308 11722 10364
rect 11658 10304 11722 10308
rect 11738 10364 11802 10368
rect 11738 10308 11742 10364
rect 11742 10308 11798 10364
rect 11798 10308 11802 10364
rect 11738 10304 11802 10308
rect 11818 10364 11882 10368
rect 11818 10308 11822 10364
rect 11822 10308 11878 10364
rect 11878 10308 11882 10364
rect 11818 10304 11882 10308
rect 11898 10364 11962 10368
rect 11898 10308 11902 10364
rect 11902 10308 11958 10364
rect 11958 10308 11962 10364
rect 11898 10304 11962 10308
rect 4010 9820 4074 9824
rect 4010 9764 4014 9820
rect 4014 9764 4070 9820
rect 4070 9764 4074 9820
rect 4010 9760 4074 9764
rect 4090 9820 4154 9824
rect 4090 9764 4094 9820
rect 4094 9764 4150 9820
rect 4150 9764 4154 9820
rect 4090 9760 4154 9764
rect 4170 9820 4234 9824
rect 4170 9764 4174 9820
rect 4174 9764 4230 9820
rect 4230 9764 4234 9820
rect 4170 9760 4234 9764
rect 4250 9820 4314 9824
rect 4250 9764 4254 9820
rect 4254 9764 4310 9820
rect 4310 9764 4314 9820
rect 4250 9760 4314 9764
rect 7069 9820 7133 9824
rect 7069 9764 7073 9820
rect 7073 9764 7129 9820
rect 7129 9764 7133 9820
rect 7069 9760 7133 9764
rect 7149 9820 7213 9824
rect 7149 9764 7153 9820
rect 7153 9764 7209 9820
rect 7209 9764 7213 9820
rect 7149 9760 7213 9764
rect 7229 9820 7293 9824
rect 7229 9764 7233 9820
rect 7233 9764 7289 9820
rect 7289 9764 7293 9820
rect 7229 9760 7293 9764
rect 7309 9820 7373 9824
rect 7309 9764 7313 9820
rect 7313 9764 7369 9820
rect 7369 9764 7373 9820
rect 7309 9760 7373 9764
rect 10128 9820 10192 9824
rect 10128 9764 10132 9820
rect 10132 9764 10188 9820
rect 10188 9764 10192 9820
rect 10128 9760 10192 9764
rect 10208 9820 10272 9824
rect 10208 9764 10212 9820
rect 10212 9764 10268 9820
rect 10268 9764 10272 9820
rect 10208 9760 10272 9764
rect 10288 9820 10352 9824
rect 10288 9764 10292 9820
rect 10292 9764 10348 9820
rect 10348 9764 10352 9820
rect 10288 9760 10352 9764
rect 10368 9820 10432 9824
rect 10368 9764 10372 9820
rect 10372 9764 10428 9820
rect 10428 9764 10432 9820
rect 10368 9760 10432 9764
rect 13187 9820 13251 9824
rect 13187 9764 13191 9820
rect 13191 9764 13247 9820
rect 13247 9764 13251 9820
rect 13187 9760 13251 9764
rect 13267 9820 13331 9824
rect 13267 9764 13271 9820
rect 13271 9764 13327 9820
rect 13327 9764 13331 9820
rect 13267 9760 13331 9764
rect 13347 9820 13411 9824
rect 13347 9764 13351 9820
rect 13351 9764 13407 9820
rect 13407 9764 13411 9820
rect 13347 9760 13411 9764
rect 13427 9820 13491 9824
rect 13427 9764 13431 9820
rect 13431 9764 13487 9820
rect 13487 9764 13491 9820
rect 13427 9760 13491 9764
rect 2481 9276 2545 9280
rect 2481 9220 2485 9276
rect 2485 9220 2541 9276
rect 2541 9220 2545 9276
rect 2481 9216 2545 9220
rect 2561 9276 2625 9280
rect 2561 9220 2565 9276
rect 2565 9220 2621 9276
rect 2621 9220 2625 9276
rect 2561 9216 2625 9220
rect 2641 9276 2705 9280
rect 2641 9220 2645 9276
rect 2645 9220 2701 9276
rect 2701 9220 2705 9276
rect 2641 9216 2705 9220
rect 2721 9276 2785 9280
rect 2721 9220 2725 9276
rect 2725 9220 2781 9276
rect 2781 9220 2785 9276
rect 2721 9216 2785 9220
rect 5540 9276 5604 9280
rect 5540 9220 5544 9276
rect 5544 9220 5600 9276
rect 5600 9220 5604 9276
rect 5540 9216 5604 9220
rect 5620 9276 5684 9280
rect 5620 9220 5624 9276
rect 5624 9220 5680 9276
rect 5680 9220 5684 9276
rect 5620 9216 5684 9220
rect 5700 9276 5764 9280
rect 5700 9220 5704 9276
rect 5704 9220 5760 9276
rect 5760 9220 5764 9276
rect 5700 9216 5764 9220
rect 5780 9276 5844 9280
rect 5780 9220 5784 9276
rect 5784 9220 5840 9276
rect 5840 9220 5844 9276
rect 5780 9216 5844 9220
rect 8599 9276 8663 9280
rect 8599 9220 8603 9276
rect 8603 9220 8659 9276
rect 8659 9220 8663 9276
rect 8599 9216 8663 9220
rect 8679 9276 8743 9280
rect 8679 9220 8683 9276
rect 8683 9220 8739 9276
rect 8739 9220 8743 9276
rect 8679 9216 8743 9220
rect 8759 9276 8823 9280
rect 8759 9220 8763 9276
rect 8763 9220 8819 9276
rect 8819 9220 8823 9276
rect 8759 9216 8823 9220
rect 8839 9276 8903 9280
rect 8839 9220 8843 9276
rect 8843 9220 8899 9276
rect 8899 9220 8903 9276
rect 8839 9216 8903 9220
rect 11658 9276 11722 9280
rect 11658 9220 11662 9276
rect 11662 9220 11718 9276
rect 11718 9220 11722 9276
rect 11658 9216 11722 9220
rect 11738 9276 11802 9280
rect 11738 9220 11742 9276
rect 11742 9220 11798 9276
rect 11798 9220 11802 9276
rect 11738 9216 11802 9220
rect 11818 9276 11882 9280
rect 11818 9220 11822 9276
rect 11822 9220 11878 9276
rect 11878 9220 11882 9276
rect 11818 9216 11882 9220
rect 11898 9276 11962 9280
rect 11898 9220 11902 9276
rect 11902 9220 11958 9276
rect 11958 9220 11962 9276
rect 11898 9216 11962 9220
rect 4010 8732 4074 8736
rect 4010 8676 4014 8732
rect 4014 8676 4070 8732
rect 4070 8676 4074 8732
rect 4010 8672 4074 8676
rect 4090 8732 4154 8736
rect 4090 8676 4094 8732
rect 4094 8676 4150 8732
rect 4150 8676 4154 8732
rect 4090 8672 4154 8676
rect 4170 8732 4234 8736
rect 4170 8676 4174 8732
rect 4174 8676 4230 8732
rect 4230 8676 4234 8732
rect 4170 8672 4234 8676
rect 4250 8732 4314 8736
rect 4250 8676 4254 8732
rect 4254 8676 4310 8732
rect 4310 8676 4314 8732
rect 4250 8672 4314 8676
rect 7069 8732 7133 8736
rect 7069 8676 7073 8732
rect 7073 8676 7129 8732
rect 7129 8676 7133 8732
rect 7069 8672 7133 8676
rect 7149 8732 7213 8736
rect 7149 8676 7153 8732
rect 7153 8676 7209 8732
rect 7209 8676 7213 8732
rect 7149 8672 7213 8676
rect 7229 8732 7293 8736
rect 7229 8676 7233 8732
rect 7233 8676 7289 8732
rect 7289 8676 7293 8732
rect 7229 8672 7293 8676
rect 7309 8732 7373 8736
rect 7309 8676 7313 8732
rect 7313 8676 7369 8732
rect 7369 8676 7373 8732
rect 7309 8672 7373 8676
rect 10128 8732 10192 8736
rect 10128 8676 10132 8732
rect 10132 8676 10188 8732
rect 10188 8676 10192 8732
rect 10128 8672 10192 8676
rect 10208 8732 10272 8736
rect 10208 8676 10212 8732
rect 10212 8676 10268 8732
rect 10268 8676 10272 8732
rect 10208 8672 10272 8676
rect 10288 8732 10352 8736
rect 10288 8676 10292 8732
rect 10292 8676 10348 8732
rect 10348 8676 10352 8732
rect 10288 8672 10352 8676
rect 10368 8732 10432 8736
rect 10368 8676 10372 8732
rect 10372 8676 10428 8732
rect 10428 8676 10432 8732
rect 10368 8672 10432 8676
rect 13187 8732 13251 8736
rect 13187 8676 13191 8732
rect 13191 8676 13247 8732
rect 13247 8676 13251 8732
rect 13187 8672 13251 8676
rect 13267 8732 13331 8736
rect 13267 8676 13271 8732
rect 13271 8676 13327 8732
rect 13327 8676 13331 8732
rect 13267 8672 13331 8676
rect 13347 8732 13411 8736
rect 13347 8676 13351 8732
rect 13351 8676 13407 8732
rect 13407 8676 13411 8732
rect 13347 8672 13411 8676
rect 13427 8732 13491 8736
rect 13427 8676 13431 8732
rect 13431 8676 13487 8732
rect 13487 8676 13491 8732
rect 13427 8672 13491 8676
rect 2481 8188 2545 8192
rect 2481 8132 2485 8188
rect 2485 8132 2541 8188
rect 2541 8132 2545 8188
rect 2481 8128 2545 8132
rect 2561 8188 2625 8192
rect 2561 8132 2565 8188
rect 2565 8132 2621 8188
rect 2621 8132 2625 8188
rect 2561 8128 2625 8132
rect 2641 8188 2705 8192
rect 2641 8132 2645 8188
rect 2645 8132 2701 8188
rect 2701 8132 2705 8188
rect 2641 8128 2705 8132
rect 2721 8188 2785 8192
rect 2721 8132 2725 8188
rect 2725 8132 2781 8188
rect 2781 8132 2785 8188
rect 2721 8128 2785 8132
rect 5540 8188 5604 8192
rect 5540 8132 5544 8188
rect 5544 8132 5600 8188
rect 5600 8132 5604 8188
rect 5540 8128 5604 8132
rect 5620 8188 5684 8192
rect 5620 8132 5624 8188
rect 5624 8132 5680 8188
rect 5680 8132 5684 8188
rect 5620 8128 5684 8132
rect 5700 8188 5764 8192
rect 5700 8132 5704 8188
rect 5704 8132 5760 8188
rect 5760 8132 5764 8188
rect 5700 8128 5764 8132
rect 5780 8188 5844 8192
rect 5780 8132 5784 8188
rect 5784 8132 5840 8188
rect 5840 8132 5844 8188
rect 5780 8128 5844 8132
rect 8599 8188 8663 8192
rect 8599 8132 8603 8188
rect 8603 8132 8659 8188
rect 8659 8132 8663 8188
rect 8599 8128 8663 8132
rect 8679 8188 8743 8192
rect 8679 8132 8683 8188
rect 8683 8132 8739 8188
rect 8739 8132 8743 8188
rect 8679 8128 8743 8132
rect 8759 8188 8823 8192
rect 8759 8132 8763 8188
rect 8763 8132 8819 8188
rect 8819 8132 8823 8188
rect 8759 8128 8823 8132
rect 8839 8188 8903 8192
rect 8839 8132 8843 8188
rect 8843 8132 8899 8188
rect 8899 8132 8903 8188
rect 8839 8128 8903 8132
rect 11658 8188 11722 8192
rect 11658 8132 11662 8188
rect 11662 8132 11718 8188
rect 11718 8132 11722 8188
rect 11658 8128 11722 8132
rect 11738 8188 11802 8192
rect 11738 8132 11742 8188
rect 11742 8132 11798 8188
rect 11798 8132 11802 8188
rect 11738 8128 11802 8132
rect 11818 8188 11882 8192
rect 11818 8132 11822 8188
rect 11822 8132 11878 8188
rect 11878 8132 11882 8188
rect 11818 8128 11882 8132
rect 11898 8188 11962 8192
rect 11898 8132 11902 8188
rect 11902 8132 11958 8188
rect 11958 8132 11962 8188
rect 11898 8128 11962 8132
rect 4010 7644 4074 7648
rect 4010 7588 4014 7644
rect 4014 7588 4070 7644
rect 4070 7588 4074 7644
rect 4010 7584 4074 7588
rect 4090 7644 4154 7648
rect 4090 7588 4094 7644
rect 4094 7588 4150 7644
rect 4150 7588 4154 7644
rect 4090 7584 4154 7588
rect 4170 7644 4234 7648
rect 4170 7588 4174 7644
rect 4174 7588 4230 7644
rect 4230 7588 4234 7644
rect 4170 7584 4234 7588
rect 4250 7644 4314 7648
rect 4250 7588 4254 7644
rect 4254 7588 4310 7644
rect 4310 7588 4314 7644
rect 4250 7584 4314 7588
rect 7069 7644 7133 7648
rect 7069 7588 7073 7644
rect 7073 7588 7129 7644
rect 7129 7588 7133 7644
rect 7069 7584 7133 7588
rect 7149 7644 7213 7648
rect 7149 7588 7153 7644
rect 7153 7588 7209 7644
rect 7209 7588 7213 7644
rect 7149 7584 7213 7588
rect 7229 7644 7293 7648
rect 7229 7588 7233 7644
rect 7233 7588 7289 7644
rect 7289 7588 7293 7644
rect 7229 7584 7293 7588
rect 7309 7644 7373 7648
rect 7309 7588 7313 7644
rect 7313 7588 7369 7644
rect 7369 7588 7373 7644
rect 7309 7584 7373 7588
rect 10128 7644 10192 7648
rect 10128 7588 10132 7644
rect 10132 7588 10188 7644
rect 10188 7588 10192 7644
rect 10128 7584 10192 7588
rect 10208 7644 10272 7648
rect 10208 7588 10212 7644
rect 10212 7588 10268 7644
rect 10268 7588 10272 7644
rect 10208 7584 10272 7588
rect 10288 7644 10352 7648
rect 10288 7588 10292 7644
rect 10292 7588 10348 7644
rect 10348 7588 10352 7644
rect 10288 7584 10352 7588
rect 10368 7644 10432 7648
rect 10368 7588 10372 7644
rect 10372 7588 10428 7644
rect 10428 7588 10432 7644
rect 10368 7584 10432 7588
rect 13187 7644 13251 7648
rect 13187 7588 13191 7644
rect 13191 7588 13247 7644
rect 13247 7588 13251 7644
rect 13187 7584 13251 7588
rect 13267 7644 13331 7648
rect 13267 7588 13271 7644
rect 13271 7588 13327 7644
rect 13327 7588 13331 7644
rect 13267 7584 13331 7588
rect 13347 7644 13411 7648
rect 13347 7588 13351 7644
rect 13351 7588 13407 7644
rect 13407 7588 13411 7644
rect 13347 7584 13411 7588
rect 13427 7644 13491 7648
rect 13427 7588 13431 7644
rect 13431 7588 13487 7644
rect 13487 7588 13491 7644
rect 13427 7584 13491 7588
rect 2481 7100 2545 7104
rect 2481 7044 2485 7100
rect 2485 7044 2541 7100
rect 2541 7044 2545 7100
rect 2481 7040 2545 7044
rect 2561 7100 2625 7104
rect 2561 7044 2565 7100
rect 2565 7044 2621 7100
rect 2621 7044 2625 7100
rect 2561 7040 2625 7044
rect 2641 7100 2705 7104
rect 2641 7044 2645 7100
rect 2645 7044 2701 7100
rect 2701 7044 2705 7100
rect 2641 7040 2705 7044
rect 2721 7100 2785 7104
rect 2721 7044 2725 7100
rect 2725 7044 2781 7100
rect 2781 7044 2785 7100
rect 2721 7040 2785 7044
rect 5540 7100 5604 7104
rect 5540 7044 5544 7100
rect 5544 7044 5600 7100
rect 5600 7044 5604 7100
rect 5540 7040 5604 7044
rect 5620 7100 5684 7104
rect 5620 7044 5624 7100
rect 5624 7044 5680 7100
rect 5680 7044 5684 7100
rect 5620 7040 5684 7044
rect 5700 7100 5764 7104
rect 5700 7044 5704 7100
rect 5704 7044 5760 7100
rect 5760 7044 5764 7100
rect 5700 7040 5764 7044
rect 5780 7100 5844 7104
rect 5780 7044 5784 7100
rect 5784 7044 5840 7100
rect 5840 7044 5844 7100
rect 5780 7040 5844 7044
rect 8599 7100 8663 7104
rect 8599 7044 8603 7100
rect 8603 7044 8659 7100
rect 8659 7044 8663 7100
rect 8599 7040 8663 7044
rect 8679 7100 8743 7104
rect 8679 7044 8683 7100
rect 8683 7044 8739 7100
rect 8739 7044 8743 7100
rect 8679 7040 8743 7044
rect 8759 7100 8823 7104
rect 8759 7044 8763 7100
rect 8763 7044 8819 7100
rect 8819 7044 8823 7100
rect 8759 7040 8823 7044
rect 8839 7100 8903 7104
rect 8839 7044 8843 7100
rect 8843 7044 8899 7100
rect 8899 7044 8903 7100
rect 8839 7040 8903 7044
rect 11658 7100 11722 7104
rect 11658 7044 11662 7100
rect 11662 7044 11718 7100
rect 11718 7044 11722 7100
rect 11658 7040 11722 7044
rect 11738 7100 11802 7104
rect 11738 7044 11742 7100
rect 11742 7044 11798 7100
rect 11798 7044 11802 7100
rect 11738 7040 11802 7044
rect 11818 7100 11882 7104
rect 11818 7044 11822 7100
rect 11822 7044 11878 7100
rect 11878 7044 11882 7100
rect 11818 7040 11882 7044
rect 11898 7100 11962 7104
rect 11898 7044 11902 7100
rect 11902 7044 11958 7100
rect 11958 7044 11962 7100
rect 11898 7040 11962 7044
rect 4010 6556 4074 6560
rect 4010 6500 4014 6556
rect 4014 6500 4070 6556
rect 4070 6500 4074 6556
rect 4010 6496 4074 6500
rect 4090 6556 4154 6560
rect 4090 6500 4094 6556
rect 4094 6500 4150 6556
rect 4150 6500 4154 6556
rect 4090 6496 4154 6500
rect 4170 6556 4234 6560
rect 4170 6500 4174 6556
rect 4174 6500 4230 6556
rect 4230 6500 4234 6556
rect 4170 6496 4234 6500
rect 4250 6556 4314 6560
rect 4250 6500 4254 6556
rect 4254 6500 4310 6556
rect 4310 6500 4314 6556
rect 4250 6496 4314 6500
rect 7069 6556 7133 6560
rect 7069 6500 7073 6556
rect 7073 6500 7129 6556
rect 7129 6500 7133 6556
rect 7069 6496 7133 6500
rect 7149 6556 7213 6560
rect 7149 6500 7153 6556
rect 7153 6500 7209 6556
rect 7209 6500 7213 6556
rect 7149 6496 7213 6500
rect 7229 6556 7293 6560
rect 7229 6500 7233 6556
rect 7233 6500 7289 6556
rect 7289 6500 7293 6556
rect 7229 6496 7293 6500
rect 7309 6556 7373 6560
rect 7309 6500 7313 6556
rect 7313 6500 7369 6556
rect 7369 6500 7373 6556
rect 7309 6496 7373 6500
rect 10128 6556 10192 6560
rect 10128 6500 10132 6556
rect 10132 6500 10188 6556
rect 10188 6500 10192 6556
rect 10128 6496 10192 6500
rect 10208 6556 10272 6560
rect 10208 6500 10212 6556
rect 10212 6500 10268 6556
rect 10268 6500 10272 6556
rect 10208 6496 10272 6500
rect 10288 6556 10352 6560
rect 10288 6500 10292 6556
rect 10292 6500 10348 6556
rect 10348 6500 10352 6556
rect 10288 6496 10352 6500
rect 10368 6556 10432 6560
rect 10368 6500 10372 6556
rect 10372 6500 10428 6556
rect 10428 6500 10432 6556
rect 10368 6496 10432 6500
rect 13187 6556 13251 6560
rect 13187 6500 13191 6556
rect 13191 6500 13247 6556
rect 13247 6500 13251 6556
rect 13187 6496 13251 6500
rect 13267 6556 13331 6560
rect 13267 6500 13271 6556
rect 13271 6500 13327 6556
rect 13327 6500 13331 6556
rect 13267 6496 13331 6500
rect 13347 6556 13411 6560
rect 13347 6500 13351 6556
rect 13351 6500 13407 6556
rect 13407 6500 13411 6556
rect 13347 6496 13411 6500
rect 13427 6556 13491 6560
rect 13427 6500 13431 6556
rect 13431 6500 13487 6556
rect 13487 6500 13491 6556
rect 13427 6496 13491 6500
rect 2481 6012 2545 6016
rect 2481 5956 2485 6012
rect 2485 5956 2541 6012
rect 2541 5956 2545 6012
rect 2481 5952 2545 5956
rect 2561 6012 2625 6016
rect 2561 5956 2565 6012
rect 2565 5956 2621 6012
rect 2621 5956 2625 6012
rect 2561 5952 2625 5956
rect 2641 6012 2705 6016
rect 2641 5956 2645 6012
rect 2645 5956 2701 6012
rect 2701 5956 2705 6012
rect 2641 5952 2705 5956
rect 2721 6012 2785 6016
rect 2721 5956 2725 6012
rect 2725 5956 2781 6012
rect 2781 5956 2785 6012
rect 2721 5952 2785 5956
rect 5540 6012 5604 6016
rect 5540 5956 5544 6012
rect 5544 5956 5600 6012
rect 5600 5956 5604 6012
rect 5540 5952 5604 5956
rect 5620 6012 5684 6016
rect 5620 5956 5624 6012
rect 5624 5956 5680 6012
rect 5680 5956 5684 6012
rect 5620 5952 5684 5956
rect 5700 6012 5764 6016
rect 5700 5956 5704 6012
rect 5704 5956 5760 6012
rect 5760 5956 5764 6012
rect 5700 5952 5764 5956
rect 5780 6012 5844 6016
rect 5780 5956 5784 6012
rect 5784 5956 5840 6012
rect 5840 5956 5844 6012
rect 5780 5952 5844 5956
rect 8599 6012 8663 6016
rect 8599 5956 8603 6012
rect 8603 5956 8659 6012
rect 8659 5956 8663 6012
rect 8599 5952 8663 5956
rect 8679 6012 8743 6016
rect 8679 5956 8683 6012
rect 8683 5956 8739 6012
rect 8739 5956 8743 6012
rect 8679 5952 8743 5956
rect 8759 6012 8823 6016
rect 8759 5956 8763 6012
rect 8763 5956 8819 6012
rect 8819 5956 8823 6012
rect 8759 5952 8823 5956
rect 8839 6012 8903 6016
rect 8839 5956 8843 6012
rect 8843 5956 8899 6012
rect 8899 5956 8903 6012
rect 8839 5952 8903 5956
rect 11658 6012 11722 6016
rect 11658 5956 11662 6012
rect 11662 5956 11718 6012
rect 11718 5956 11722 6012
rect 11658 5952 11722 5956
rect 11738 6012 11802 6016
rect 11738 5956 11742 6012
rect 11742 5956 11798 6012
rect 11798 5956 11802 6012
rect 11738 5952 11802 5956
rect 11818 6012 11882 6016
rect 11818 5956 11822 6012
rect 11822 5956 11878 6012
rect 11878 5956 11882 6012
rect 11818 5952 11882 5956
rect 11898 6012 11962 6016
rect 11898 5956 11902 6012
rect 11902 5956 11958 6012
rect 11958 5956 11962 6012
rect 11898 5952 11962 5956
rect 4010 5468 4074 5472
rect 4010 5412 4014 5468
rect 4014 5412 4070 5468
rect 4070 5412 4074 5468
rect 4010 5408 4074 5412
rect 4090 5468 4154 5472
rect 4090 5412 4094 5468
rect 4094 5412 4150 5468
rect 4150 5412 4154 5468
rect 4090 5408 4154 5412
rect 4170 5468 4234 5472
rect 4170 5412 4174 5468
rect 4174 5412 4230 5468
rect 4230 5412 4234 5468
rect 4170 5408 4234 5412
rect 4250 5468 4314 5472
rect 4250 5412 4254 5468
rect 4254 5412 4310 5468
rect 4310 5412 4314 5468
rect 4250 5408 4314 5412
rect 7069 5468 7133 5472
rect 7069 5412 7073 5468
rect 7073 5412 7129 5468
rect 7129 5412 7133 5468
rect 7069 5408 7133 5412
rect 7149 5468 7213 5472
rect 7149 5412 7153 5468
rect 7153 5412 7209 5468
rect 7209 5412 7213 5468
rect 7149 5408 7213 5412
rect 7229 5468 7293 5472
rect 7229 5412 7233 5468
rect 7233 5412 7289 5468
rect 7289 5412 7293 5468
rect 7229 5408 7293 5412
rect 7309 5468 7373 5472
rect 7309 5412 7313 5468
rect 7313 5412 7369 5468
rect 7369 5412 7373 5468
rect 7309 5408 7373 5412
rect 10128 5468 10192 5472
rect 10128 5412 10132 5468
rect 10132 5412 10188 5468
rect 10188 5412 10192 5468
rect 10128 5408 10192 5412
rect 10208 5468 10272 5472
rect 10208 5412 10212 5468
rect 10212 5412 10268 5468
rect 10268 5412 10272 5468
rect 10208 5408 10272 5412
rect 10288 5468 10352 5472
rect 10288 5412 10292 5468
rect 10292 5412 10348 5468
rect 10348 5412 10352 5468
rect 10288 5408 10352 5412
rect 10368 5468 10432 5472
rect 10368 5412 10372 5468
rect 10372 5412 10428 5468
rect 10428 5412 10432 5468
rect 10368 5408 10432 5412
rect 13187 5468 13251 5472
rect 13187 5412 13191 5468
rect 13191 5412 13247 5468
rect 13247 5412 13251 5468
rect 13187 5408 13251 5412
rect 13267 5468 13331 5472
rect 13267 5412 13271 5468
rect 13271 5412 13327 5468
rect 13327 5412 13331 5468
rect 13267 5408 13331 5412
rect 13347 5468 13411 5472
rect 13347 5412 13351 5468
rect 13351 5412 13407 5468
rect 13407 5412 13411 5468
rect 13347 5408 13411 5412
rect 13427 5468 13491 5472
rect 13427 5412 13431 5468
rect 13431 5412 13487 5468
rect 13487 5412 13491 5468
rect 13427 5408 13491 5412
rect 2481 4924 2545 4928
rect 2481 4868 2485 4924
rect 2485 4868 2541 4924
rect 2541 4868 2545 4924
rect 2481 4864 2545 4868
rect 2561 4924 2625 4928
rect 2561 4868 2565 4924
rect 2565 4868 2621 4924
rect 2621 4868 2625 4924
rect 2561 4864 2625 4868
rect 2641 4924 2705 4928
rect 2641 4868 2645 4924
rect 2645 4868 2701 4924
rect 2701 4868 2705 4924
rect 2641 4864 2705 4868
rect 2721 4924 2785 4928
rect 2721 4868 2725 4924
rect 2725 4868 2781 4924
rect 2781 4868 2785 4924
rect 2721 4864 2785 4868
rect 5540 4924 5604 4928
rect 5540 4868 5544 4924
rect 5544 4868 5600 4924
rect 5600 4868 5604 4924
rect 5540 4864 5604 4868
rect 5620 4924 5684 4928
rect 5620 4868 5624 4924
rect 5624 4868 5680 4924
rect 5680 4868 5684 4924
rect 5620 4864 5684 4868
rect 5700 4924 5764 4928
rect 5700 4868 5704 4924
rect 5704 4868 5760 4924
rect 5760 4868 5764 4924
rect 5700 4864 5764 4868
rect 5780 4924 5844 4928
rect 5780 4868 5784 4924
rect 5784 4868 5840 4924
rect 5840 4868 5844 4924
rect 5780 4864 5844 4868
rect 8599 4924 8663 4928
rect 8599 4868 8603 4924
rect 8603 4868 8659 4924
rect 8659 4868 8663 4924
rect 8599 4864 8663 4868
rect 8679 4924 8743 4928
rect 8679 4868 8683 4924
rect 8683 4868 8739 4924
rect 8739 4868 8743 4924
rect 8679 4864 8743 4868
rect 8759 4924 8823 4928
rect 8759 4868 8763 4924
rect 8763 4868 8819 4924
rect 8819 4868 8823 4924
rect 8759 4864 8823 4868
rect 8839 4924 8903 4928
rect 8839 4868 8843 4924
rect 8843 4868 8899 4924
rect 8899 4868 8903 4924
rect 8839 4864 8903 4868
rect 11658 4924 11722 4928
rect 11658 4868 11662 4924
rect 11662 4868 11718 4924
rect 11718 4868 11722 4924
rect 11658 4864 11722 4868
rect 11738 4924 11802 4928
rect 11738 4868 11742 4924
rect 11742 4868 11798 4924
rect 11798 4868 11802 4924
rect 11738 4864 11802 4868
rect 11818 4924 11882 4928
rect 11818 4868 11822 4924
rect 11822 4868 11878 4924
rect 11878 4868 11882 4924
rect 11818 4864 11882 4868
rect 11898 4924 11962 4928
rect 11898 4868 11902 4924
rect 11902 4868 11958 4924
rect 11958 4868 11962 4924
rect 11898 4864 11962 4868
rect 4010 4380 4074 4384
rect 4010 4324 4014 4380
rect 4014 4324 4070 4380
rect 4070 4324 4074 4380
rect 4010 4320 4074 4324
rect 4090 4380 4154 4384
rect 4090 4324 4094 4380
rect 4094 4324 4150 4380
rect 4150 4324 4154 4380
rect 4090 4320 4154 4324
rect 4170 4380 4234 4384
rect 4170 4324 4174 4380
rect 4174 4324 4230 4380
rect 4230 4324 4234 4380
rect 4170 4320 4234 4324
rect 4250 4380 4314 4384
rect 4250 4324 4254 4380
rect 4254 4324 4310 4380
rect 4310 4324 4314 4380
rect 4250 4320 4314 4324
rect 7069 4380 7133 4384
rect 7069 4324 7073 4380
rect 7073 4324 7129 4380
rect 7129 4324 7133 4380
rect 7069 4320 7133 4324
rect 7149 4380 7213 4384
rect 7149 4324 7153 4380
rect 7153 4324 7209 4380
rect 7209 4324 7213 4380
rect 7149 4320 7213 4324
rect 7229 4380 7293 4384
rect 7229 4324 7233 4380
rect 7233 4324 7289 4380
rect 7289 4324 7293 4380
rect 7229 4320 7293 4324
rect 7309 4380 7373 4384
rect 7309 4324 7313 4380
rect 7313 4324 7369 4380
rect 7369 4324 7373 4380
rect 7309 4320 7373 4324
rect 10128 4380 10192 4384
rect 10128 4324 10132 4380
rect 10132 4324 10188 4380
rect 10188 4324 10192 4380
rect 10128 4320 10192 4324
rect 10208 4380 10272 4384
rect 10208 4324 10212 4380
rect 10212 4324 10268 4380
rect 10268 4324 10272 4380
rect 10208 4320 10272 4324
rect 10288 4380 10352 4384
rect 10288 4324 10292 4380
rect 10292 4324 10348 4380
rect 10348 4324 10352 4380
rect 10288 4320 10352 4324
rect 10368 4380 10432 4384
rect 10368 4324 10372 4380
rect 10372 4324 10428 4380
rect 10428 4324 10432 4380
rect 10368 4320 10432 4324
rect 13187 4380 13251 4384
rect 13187 4324 13191 4380
rect 13191 4324 13247 4380
rect 13247 4324 13251 4380
rect 13187 4320 13251 4324
rect 13267 4380 13331 4384
rect 13267 4324 13271 4380
rect 13271 4324 13327 4380
rect 13327 4324 13331 4380
rect 13267 4320 13331 4324
rect 13347 4380 13411 4384
rect 13347 4324 13351 4380
rect 13351 4324 13407 4380
rect 13407 4324 13411 4380
rect 13347 4320 13411 4324
rect 13427 4380 13491 4384
rect 13427 4324 13431 4380
rect 13431 4324 13487 4380
rect 13487 4324 13491 4380
rect 13427 4320 13491 4324
rect 2481 3836 2545 3840
rect 2481 3780 2485 3836
rect 2485 3780 2541 3836
rect 2541 3780 2545 3836
rect 2481 3776 2545 3780
rect 2561 3836 2625 3840
rect 2561 3780 2565 3836
rect 2565 3780 2621 3836
rect 2621 3780 2625 3836
rect 2561 3776 2625 3780
rect 2641 3836 2705 3840
rect 2641 3780 2645 3836
rect 2645 3780 2701 3836
rect 2701 3780 2705 3836
rect 2641 3776 2705 3780
rect 2721 3836 2785 3840
rect 2721 3780 2725 3836
rect 2725 3780 2781 3836
rect 2781 3780 2785 3836
rect 2721 3776 2785 3780
rect 5540 3836 5604 3840
rect 5540 3780 5544 3836
rect 5544 3780 5600 3836
rect 5600 3780 5604 3836
rect 5540 3776 5604 3780
rect 5620 3836 5684 3840
rect 5620 3780 5624 3836
rect 5624 3780 5680 3836
rect 5680 3780 5684 3836
rect 5620 3776 5684 3780
rect 5700 3836 5764 3840
rect 5700 3780 5704 3836
rect 5704 3780 5760 3836
rect 5760 3780 5764 3836
rect 5700 3776 5764 3780
rect 5780 3836 5844 3840
rect 5780 3780 5784 3836
rect 5784 3780 5840 3836
rect 5840 3780 5844 3836
rect 5780 3776 5844 3780
rect 8599 3836 8663 3840
rect 8599 3780 8603 3836
rect 8603 3780 8659 3836
rect 8659 3780 8663 3836
rect 8599 3776 8663 3780
rect 8679 3836 8743 3840
rect 8679 3780 8683 3836
rect 8683 3780 8739 3836
rect 8739 3780 8743 3836
rect 8679 3776 8743 3780
rect 8759 3836 8823 3840
rect 8759 3780 8763 3836
rect 8763 3780 8819 3836
rect 8819 3780 8823 3836
rect 8759 3776 8823 3780
rect 8839 3836 8903 3840
rect 8839 3780 8843 3836
rect 8843 3780 8899 3836
rect 8899 3780 8903 3836
rect 8839 3776 8903 3780
rect 11658 3836 11722 3840
rect 11658 3780 11662 3836
rect 11662 3780 11718 3836
rect 11718 3780 11722 3836
rect 11658 3776 11722 3780
rect 11738 3836 11802 3840
rect 11738 3780 11742 3836
rect 11742 3780 11798 3836
rect 11798 3780 11802 3836
rect 11738 3776 11802 3780
rect 11818 3836 11882 3840
rect 11818 3780 11822 3836
rect 11822 3780 11878 3836
rect 11878 3780 11882 3836
rect 11818 3776 11882 3780
rect 11898 3836 11962 3840
rect 11898 3780 11902 3836
rect 11902 3780 11958 3836
rect 11958 3780 11962 3836
rect 11898 3776 11962 3780
rect 4010 3292 4074 3296
rect 4010 3236 4014 3292
rect 4014 3236 4070 3292
rect 4070 3236 4074 3292
rect 4010 3232 4074 3236
rect 4090 3292 4154 3296
rect 4090 3236 4094 3292
rect 4094 3236 4150 3292
rect 4150 3236 4154 3292
rect 4090 3232 4154 3236
rect 4170 3292 4234 3296
rect 4170 3236 4174 3292
rect 4174 3236 4230 3292
rect 4230 3236 4234 3292
rect 4170 3232 4234 3236
rect 4250 3292 4314 3296
rect 4250 3236 4254 3292
rect 4254 3236 4310 3292
rect 4310 3236 4314 3292
rect 4250 3232 4314 3236
rect 7069 3292 7133 3296
rect 7069 3236 7073 3292
rect 7073 3236 7129 3292
rect 7129 3236 7133 3292
rect 7069 3232 7133 3236
rect 7149 3292 7213 3296
rect 7149 3236 7153 3292
rect 7153 3236 7209 3292
rect 7209 3236 7213 3292
rect 7149 3232 7213 3236
rect 7229 3292 7293 3296
rect 7229 3236 7233 3292
rect 7233 3236 7289 3292
rect 7289 3236 7293 3292
rect 7229 3232 7293 3236
rect 7309 3292 7373 3296
rect 7309 3236 7313 3292
rect 7313 3236 7369 3292
rect 7369 3236 7373 3292
rect 7309 3232 7373 3236
rect 10128 3292 10192 3296
rect 10128 3236 10132 3292
rect 10132 3236 10188 3292
rect 10188 3236 10192 3292
rect 10128 3232 10192 3236
rect 10208 3292 10272 3296
rect 10208 3236 10212 3292
rect 10212 3236 10268 3292
rect 10268 3236 10272 3292
rect 10208 3232 10272 3236
rect 10288 3292 10352 3296
rect 10288 3236 10292 3292
rect 10292 3236 10348 3292
rect 10348 3236 10352 3292
rect 10288 3232 10352 3236
rect 10368 3292 10432 3296
rect 10368 3236 10372 3292
rect 10372 3236 10428 3292
rect 10428 3236 10432 3292
rect 10368 3232 10432 3236
rect 13187 3292 13251 3296
rect 13187 3236 13191 3292
rect 13191 3236 13247 3292
rect 13247 3236 13251 3292
rect 13187 3232 13251 3236
rect 13267 3292 13331 3296
rect 13267 3236 13271 3292
rect 13271 3236 13327 3292
rect 13327 3236 13331 3292
rect 13267 3232 13331 3236
rect 13347 3292 13411 3296
rect 13347 3236 13351 3292
rect 13351 3236 13407 3292
rect 13407 3236 13411 3292
rect 13347 3232 13411 3236
rect 13427 3292 13491 3296
rect 13427 3236 13431 3292
rect 13431 3236 13487 3292
rect 13487 3236 13491 3292
rect 13427 3232 13491 3236
rect 2481 2748 2545 2752
rect 2481 2692 2485 2748
rect 2485 2692 2541 2748
rect 2541 2692 2545 2748
rect 2481 2688 2545 2692
rect 2561 2748 2625 2752
rect 2561 2692 2565 2748
rect 2565 2692 2621 2748
rect 2621 2692 2625 2748
rect 2561 2688 2625 2692
rect 2641 2748 2705 2752
rect 2641 2692 2645 2748
rect 2645 2692 2701 2748
rect 2701 2692 2705 2748
rect 2641 2688 2705 2692
rect 2721 2748 2785 2752
rect 2721 2692 2725 2748
rect 2725 2692 2781 2748
rect 2781 2692 2785 2748
rect 2721 2688 2785 2692
rect 5540 2748 5604 2752
rect 5540 2692 5544 2748
rect 5544 2692 5600 2748
rect 5600 2692 5604 2748
rect 5540 2688 5604 2692
rect 5620 2748 5684 2752
rect 5620 2692 5624 2748
rect 5624 2692 5680 2748
rect 5680 2692 5684 2748
rect 5620 2688 5684 2692
rect 5700 2748 5764 2752
rect 5700 2692 5704 2748
rect 5704 2692 5760 2748
rect 5760 2692 5764 2748
rect 5700 2688 5764 2692
rect 5780 2748 5844 2752
rect 5780 2692 5784 2748
rect 5784 2692 5840 2748
rect 5840 2692 5844 2748
rect 5780 2688 5844 2692
rect 8599 2748 8663 2752
rect 8599 2692 8603 2748
rect 8603 2692 8659 2748
rect 8659 2692 8663 2748
rect 8599 2688 8663 2692
rect 8679 2748 8743 2752
rect 8679 2692 8683 2748
rect 8683 2692 8739 2748
rect 8739 2692 8743 2748
rect 8679 2688 8743 2692
rect 8759 2748 8823 2752
rect 8759 2692 8763 2748
rect 8763 2692 8819 2748
rect 8819 2692 8823 2748
rect 8759 2688 8823 2692
rect 8839 2748 8903 2752
rect 8839 2692 8843 2748
rect 8843 2692 8899 2748
rect 8899 2692 8903 2748
rect 8839 2688 8903 2692
rect 11658 2748 11722 2752
rect 11658 2692 11662 2748
rect 11662 2692 11718 2748
rect 11718 2692 11722 2748
rect 11658 2688 11722 2692
rect 11738 2748 11802 2752
rect 11738 2692 11742 2748
rect 11742 2692 11798 2748
rect 11798 2692 11802 2748
rect 11738 2688 11802 2692
rect 11818 2748 11882 2752
rect 11818 2692 11822 2748
rect 11822 2692 11878 2748
rect 11878 2692 11882 2748
rect 11818 2688 11882 2692
rect 11898 2748 11962 2752
rect 11898 2692 11902 2748
rect 11902 2692 11958 2748
rect 11958 2692 11962 2748
rect 11898 2688 11962 2692
rect 4010 2204 4074 2208
rect 4010 2148 4014 2204
rect 4014 2148 4070 2204
rect 4070 2148 4074 2204
rect 4010 2144 4074 2148
rect 4090 2204 4154 2208
rect 4090 2148 4094 2204
rect 4094 2148 4150 2204
rect 4150 2148 4154 2204
rect 4090 2144 4154 2148
rect 4170 2204 4234 2208
rect 4170 2148 4174 2204
rect 4174 2148 4230 2204
rect 4230 2148 4234 2204
rect 4170 2144 4234 2148
rect 4250 2204 4314 2208
rect 4250 2148 4254 2204
rect 4254 2148 4310 2204
rect 4310 2148 4314 2204
rect 4250 2144 4314 2148
rect 7069 2204 7133 2208
rect 7069 2148 7073 2204
rect 7073 2148 7129 2204
rect 7129 2148 7133 2204
rect 7069 2144 7133 2148
rect 7149 2204 7213 2208
rect 7149 2148 7153 2204
rect 7153 2148 7209 2204
rect 7209 2148 7213 2204
rect 7149 2144 7213 2148
rect 7229 2204 7293 2208
rect 7229 2148 7233 2204
rect 7233 2148 7289 2204
rect 7289 2148 7293 2204
rect 7229 2144 7293 2148
rect 7309 2204 7373 2208
rect 7309 2148 7313 2204
rect 7313 2148 7369 2204
rect 7369 2148 7373 2204
rect 7309 2144 7373 2148
rect 10128 2204 10192 2208
rect 10128 2148 10132 2204
rect 10132 2148 10188 2204
rect 10188 2148 10192 2204
rect 10128 2144 10192 2148
rect 10208 2204 10272 2208
rect 10208 2148 10212 2204
rect 10212 2148 10268 2204
rect 10268 2148 10272 2204
rect 10208 2144 10272 2148
rect 10288 2204 10352 2208
rect 10288 2148 10292 2204
rect 10292 2148 10348 2204
rect 10348 2148 10352 2204
rect 10288 2144 10352 2148
rect 10368 2204 10432 2208
rect 10368 2148 10372 2204
rect 10372 2148 10428 2204
rect 10428 2148 10432 2204
rect 10368 2144 10432 2148
rect 13187 2204 13251 2208
rect 13187 2148 13191 2204
rect 13191 2148 13247 2204
rect 13247 2148 13251 2204
rect 13187 2144 13251 2148
rect 13267 2204 13331 2208
rect 13267 2148 13271 2204
rect 13271 2148 13327 2204
rect 13327 2148 13331 2204
rect 13267 2144 13331 2148
rect 13347 2204 13411 2208
rect 13347 2148 13351 2204
rect 13351 2148 13407 2204
rect 13407 2148 13411 2204
rect 13347 2144 13411 2148
rect 13427 2204 13491 2208
rect 13427 2148 13431 2204
rect 13431 2148 13487 2204
rect 13487 2148 13491 2204
rect 13427 2144 13491 2148
<< metal4 >>
rect 2473 13632 2793 14192
rect 2473 13568 2481 13632
rect 2545 13568 2561 13632
rect 2625 13568 2641 13632
rect 2705 13568 2721 13632
rect 2785 13568 2793 13632
rect 2473 12544 2793 13568
rect 2473 12480 2481 12544
rect 2545 12480 2561 12544
rect 2625 12480 2641 12544
rect 2705 12480 2721 12544
rect 2785 12480 2793 12544
rect 2473 11456 2793 12480
rect 2473 11392 2481 11456
rect 2545 11392 2561 11456
rect 2625 11392 2641 11456
rect 2705 11392 2721 11456
rect 2785 11392 2793 11456
rect 2473 10368 2793 11392
rect 2473 10304 2481 10368
rect 2545 10304 2561 10368
rect 2625 10304 2641 10368
rect 2705 10304 2721 10368
rect 2785 10304 2793 10368
rect 2473 9280 2793 10304
rect 2473 9216 2481 9280
rect 2545 9216 2561 9280
rect 2625 9216 2641 9280
rect 2705 9216 2721 9280
rect 2785 9216 2793 9280
rect 2473 8192 2793 9216
rect 2473 8128 2481 8192
rect 2545 8128 2561 8192
rect 2625 8128 2641 8192
rect 2705 8128 2721 8192
rect 2785 8128 2793 8192
rect 2473 7104 2793 8128
rect 2473 7040 2481 7104
rect 2545 7040 2561 7104
rect 2625 7040 2641 7104
rect 2705 7040 2721 7104
rect 2785 7040 2793 7104
rect 2473 6016 2793 7040
rect 2473 5952 2481 6016
rect 2545 5952 2561 6016
rect 2625 5952 2641 6016
rect 2705 5952 2721 6016
rect 2785 5952 2793 6016
rect 2473 4928 2793 5952
rect 2473 4864 2481 4928
rect 2545 4864 2561 4928
rect 2625 4864 2641 4928
rect 2705 4864 2721 4928
rect 2785 4864 2793 4928
rect 2473 3840 2793 4864
rect 2473 3776 2481 3840
rect 2545 3776 2561 3840
rect 2625 3776 2641 3840
rect 2705 3776 2721 3840
rect 2785 3776 2793 3840
rect 2473 2752 2793 3776
rect 2473 2688 2481 2752
rect 2545 2688 2561 2752
rect 2625 2688 2641 2752
rect 2705 2688 2721 2752
rect 2785 2688 2793 2752
rect 2473 2128 2793 2688
rect 4002 14176 4322 14192
rect 4002 14112 4010 14176
rect 4074 14112 4090 14176
rect 4154 14112 4170 14176
rect 4234 14112 4250 14176
rect 4314 14112 4322 14176
rect 4002 13088 4322 14112
rect 4002 13024 4010 13088
rect 4074 13024 4090 13088
rect 4154 13024 4170 13088
rect 4234 13024 4250 13088
rect 4314 13024 4322 13088
rect 4002 12000 4322 13024
rect 4002 11936 4010 12000
rect 4074 11936 4090 12000
rect 4154 11936 4170 12000
rect 4234 11936 4250 12000
rect 4314 11936 4322 12000
rect 4002 10912 4322 11936
rect 4002 10848 4010 10912
rect 4074 10848 4090 10912
rect 4154 10848 4170 10912
rect 4234 10848 4250 10912
rect 4314 10848 4322 10912
rect 4002 9824 4322 10848
rect 4002 9760 4010 9824
rect 4074 9760 4090 9824
rect 4154 9760 4170 9824
rect 4234 9760 4250 9824
rect 4314 9760 4322 9824
rect 4002 8736 4322 9760
rect 4002 8672 4010 8736
rect 4074 8672 4090 8736
rect 4154 8672 4170 8736
rect 4234 8672 4250 8736
rect 4314 8672 4322 8736
rect 4002 7648 4322 8672
rect 4002 7584 4010 7648
rect 4074 7584 4090 7648
rect 4154 7584 4170 7648
rect 4234 7584 4250 7648
rect 4314 7584 4322 7648
rect 4002 6560 4322 7584
rect 4002 6496 4010 6560
rect 4074 6496 4090 6560
rect 4154 6496 4170 6560
rect 4234 6496 4250 6560
rect 4314 6496 4322 6560
rect 4002 5472 4322 6496
rect 4002 5408 4010 5472
rect 4074 5408 4090 5472
rect 4154 5408 4170 5472
rect 4234 5408 4250 5472
rect 4314 5408 4322 5472
rect 4002 4384 4322 5408
rect 4002 4320 4010 4384
rect 4074 4320 4090 4384
rect 4154 4320 4170 4384
rect 4234 4320 4250 4384
rect 4314 4320 4322 4384
rect 4002 3296 4322 4320
rect 4002 3232 4010 3296
rect 4074 3232 4090 3296
rect 4154 3232 4170 3296
rect 4234 3232 4250 3296
rect 4314 3232 4322 3296
rect 4002 2208 4322 3232
rect 4002 2144 4010 2208
rect 4074 2144 4090 2208
rect 4154 2144 4170 2208
rect 4234 2144 4250 2208
rect 4314 2144 4322 2208
rect 4002 2128 4322 2144
rect 5532 13632 5852 14192
rect 5532 13568 5540 13632
rect 5604 13568 5620 13632
rect 5684 13568 5700 13632
rect 5764 13568 5780 13632
rect 5844 13568 5852 13632
rect 5532 12544 5852 13568
rect 5532 12480 5540 12544
rect 5604 12480 5620 12544
rect 5684 12480 5700 12544
rect 5764 12480 5780 12544
rect 5844 12480 5852 12544
rect 5532 11456 5852 12480
rect 5532 11392 5540 11456
rect 5604 11392 5620 11456
rect 5684 11392 5700 11456
rect 5764 11392 5780 11456
rect 5844 11392 5852 11456
rect 5532 10368 5852 11392
rect 5532 10304 5540 10368
rect 5604 10304 5620 10368
rect 5684 10304 5700 10368
rect 5764 10304 5780 10368
rect 5844 10304 5852 10368
rect 5532 9280 5852 10304
rect 5532 9216 5540 9280
rect 5604 9216 5620 9280
rect 5684 9216 5700 9280
rect 5764 9216 5780 9280
rect 5844 9216 5852 9280
rect 5532 8192 5852 9216
rect 5532 8128 5540 8192
rect 5604 8128 5620 8192
rect 5684 8128 5700 8192
rect 5764 8128 5780 8192
rect 5844 8128 5852 8192
rect 5532 7104 5852 8128
rect 5532 7040 5540 7104
rect 5604 7040 5620 7104
rect 5684 7040 5700 7104
rect 5764 7040 5780 7104
rect 5844 7040 5852 7104
rect 5532 6016 5852 7040
rect 5532 5952 5540 6016
rect 5604 5952 5620 6016
rect 5684 5952 5700 6016
rect 5764 5952 5780 6016
rect 5844 5952 5852 6016
rect 5532 4928 5852 5952
rect 5532 4864 5540 4928
rect 5604 4864 5620 4928
rect 5684 4864 5700 4928
rect 5764 4864 5780 4928
rect 5844 4864 5852 4928
rect 5532 3840 5852 4864
rect 5532 3776 5540 3840
rect 5604 3776 5620 3840
rect 5684 3776 5700 3840
rect 5764 3776 5780 3840
rect 5844 3776 5852 3840
rect 5532 2752 5852 3776
rect 5532 2688 5540 2752
rect 5604 2688 5620 2752
rect 5684 2688 5700 2752
rect 5764 2688 5780 2752
rect 5844 2688 5852 2752
rect 5532 2128 5852 2688
rect 7061 14176 7381 14192
rect 7061 14112 7069 14176
rect 7133 14112 7149 14176
rect 7213 14112 7229 14176
rect 7293 14112 7309 14176
rect 7373 14112 7381 14176
rect 7061 13088 7381 14112
rect 7061 13024 7069 13088
rect 7133 13024 7149 13088
rect 7213 13024 7229 13088
rect 7293 13024 7309 13088
rect 7373 13024 7381 13088
rect 7061 12000 7381 13024
rect 7061 11936 7069 12000
rect 7133 11936 7149 12000
rect 7213 11936 7229 12000
rect 7293 11936 7309 12000
rect 7373 11936 7381 12000
rect 7061 10912 7381 11936
rect 7061 10848 7069 10912
rect 7133 10848 7149 10912
rect 7213 10848 7229 10912
rect 7293 10848 7309 10912
rect 7373 10848 7381 10912
rect 7061 9824 7381 10848
rect 7061 9760 7069 9824
rect 7133 9760 7149 9824
rect 7213 9760 7229 9824
rect 7293 9760 7309 9824
rect 7373 9760 7381 9824
rect 7061 8736 7381 9760
rect 7061 8672 7069 8736
rect 7133 8672 7149 8736
rect 7213 8672 7229 8736
rect 7293 8672 7309 8736
rect 7373 8672 7381 8736
rect 7061 7648 7381 8672
rect 7061 7584 7069 7648
rect 7133 7584 7149 7648
rect 7213 7584 7229 7648
rect 7293 7584 7309 7648
rect 7373 7584 7381 7648
rect 7061 6560 7381 7584
rect 7061 6496 7069 6560
rect 7133 6496 7149 6560
rect 7213 6496 7229 6560
rect 7293 6496 7309 6560
rect 7373 6496 7381 6560
rect 7061 5472 7381 6496
rect 7061 5408 7069 5472
rect 7133 5408 7149 5472
rect 7213 5408 7229 5472
rect 7293 5408 7309 5472
rect 7373 5408 7381 5472
rect 7061 4384 7381 5408
rect 7061 4320 7069 4384
rect 7133 4320 7149 4384
rect 7213 4320 7229 4384
rect 7293 4320 7309 4384
rect 7373 4320 7381 4384
rect 7061 3296 7381 4320
rect 7061 3232 7069 3296
rect 7133 3232 7149 3296
rect 7213 3232 7229 3296
rect 7293 3232 7309 3296
rect 7373 3232 7381 3296
rect 7061 2208 7381 3232
rect 7061 2144 7069 2208
rect 7133 2144 7149 2208
rect 7213 2144 7229 2208
rect 7293 2144 7309 2208
rect 7373 2144 7381 2208
rect 7061 2128 7381 2144
rect 8591 13632 8911 14192
rect 8591 13568 8599 13632
rect 8663 13568 8679 13632
rect 8743 13568 8759 13632
rect 8823 13568 8839 13632
rect 8903 13568 8911 13632
rect 8591 12544 8911 13568
rect 8591 12480 8599 12544
rect 8663 12480 8679 12544
rect 8743 12480 8759 12544
rect 8823 12480 8839 12544
rect 8903 12480 8911 12544
rect 8591 11456 8911 12480
rect 8591 11392 8599 11456
rect 8663 11392 8679 11456
rect 8743 11392 8759 11456
rect 8823 11392 8839 11456
rect 8903 11392 8911 11456
rect 8591 10368 8911 11392
rect 8591 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8911 10368
rect 8591 9280 8911 10304
rect 8591 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8911 9280
rect 8591 8192 8911 9216
rect 8591 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8911 8192
rect 8591 7104 8911 8128
rect 8591 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8911 7104
rect 8591 6016 8911 7040
rect 8591 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8911 6016
rect 8591 4928 8911 5952
rect 8591 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8911 4928
rect 8591 3840 8911 4864
rect 8591 3776 8599 3840
rect 8663 3776 8679 3840
rect 8743 3776 8759 3840
rect 8823 3776 8839 3840
rect 8903 3776 8911 3840
rect 8591 2752 8911 3776
rect 8591 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8911 2752
rect 8591 2128 8911 2688
rect 10120 14176 10440 14192
rect 10120 14112 10128 14176
rect 10192 14112 10208 14176
rect 10272 14112 10288 14176
rect 10352 14112 10368 14176
rect 10432 14112 10440 14176
rect 10120 13088 10440 14112
rect 10120 13024 10128 13088
rect 10192 13024 10208 13088
rect 10272 13024 10288 13088
rect 10352 13024 10368 13088
rect 10432 13024 10440 13088
rect 10120 12000 10440 13024
rect 10120 11936 10128 12000
rect 10192 11936 10208 12000
rect 10272 11936 10288 12000
rect 10352 11936 10368 12000
rect 10432 11936 10440 12000
rect 10120 10912 10440 11936
rect 10120 10848 10128 10912
rect 10192 10848 10208 10912
rect 10272 10848 10288 10912
rect 10352 10848 10368 10912
rect 10432 10848 10440 10912
rect 10120 9824 10440 10848
rect 10120 9760 10128 9824
rect 10192 9760 10208 9824
rect 10272 9760 10288 9824
rect 10352 9760 10368 9824
rect 10432 9760 10440 9824
rect 10120 8736 10440 9760
rect 10120 8672 10128 8736
rect 10192 8672 10208 8736
rect 10272 8672 10288 8736
rect 10352 8672 10368 8736
rect 10432 8672 10440 8736
rect 10120 7648 10440 8672
rect 10120 7584 10128 7648
rect 10192 7584 10208 7648
rect 10272 7584 10288 7648
rect 10352 7584 10368 7648
rect 10432 7584 10440 7648
rect 10120 6560 10440 7584
rect 10120 6496 10128 6560
rect 10192 6496 10208 6560
rect 10272 6496 10288 6560
rect 10352 6496 10368 6560
rect 10432 6496 10440 6560
rect 10120 5472 10440 6496
rect 10120 5408 10128 5472
rect 10192 5408 10208 5472
rect 10272 5408 10288 5472
rect 10352 5408 10368 5472
rect 10432 5408 10440 5472
rect 10120 4384 10440 5408
rect 10120 4320 10128 4384
rect 10192 4320 10208 4384
rect 10272 4320 10288 4384
rect 10352 4320 10368 4384
rect 10432 4320 10440 4384
rect 10120 3296 10440 4320
rect 10120 3232 10128 3296
rect 10192 3232 10208 3296
rect 10272 3232 10288 3296
rect 10352 3232 10368 3296
rect 10432 3232 10440 3296
rect 10120 2208 10440 3232
rect 10120 2144 10128 2208
rect 10192 2144 10208 2208
rect 10272 2144 10288 2208
rect 10352 2144 10368 2208
rect 10432 2144 10440 2208
rect 10120 2128 10440 2144
rect 11650 13632 11970 14192
rect 11650 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11898 13632
rect 11962 13568 11970 13632
rect 11650 12544 11970 13568
rect 11650 12480 11658 12544
rect 11722 12480 11738 12544
rect 11802 12480 11818 12544
rect 11882 12480 11898 12544
rect 11962 12480 11970 12544
rect 11650 11456 11970 12480
rect 11650 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11898 11456
rect 11962 11392 11970 11456
rect 11650 10368 11970 11392
rect 11650 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11898 10368
rect 11962 10304 11970 10368
rect 11650 9280 11970 10304
rect 11650 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11898 9280
rect 11962 9216 11970 9280
rect 11650 8192 11970 9216
rect 11650 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11898 8192
rect 11962 8128 11970 8192
rect 11650 7104 11970 8128
rect 11650 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11898 7104
rect 11962 7040 11970 7104
rect 11650 6016 11970 7040
rect 11650 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11898 6016
rect 11962 5952 11970 6016
rect 11650 4928 11970 5952
rect 11650 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11898 4928
rect 11962 4864 11970 4928
rect 11650 3840 11970 4864
rect 11650 3776 11658 3840
rect 11722 3776 11738 3840
rect 11802 3776 11818 3840
rect 11882 3776 11898 3840
rect 11962 3776 11970 3840
rect 11650 2752 11970 3776
rect 11650 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11898 2752
rect 11962 2688 11970 2752
rect 11650 2128 11970 2688
rect 13179 14176 13499 14192
rect 13179 14112 13187 14176
rect 13251 14112 13267 14176
rect 13331 14112 13347 14176
rect 13411 14112 13427 14176
rect 13491 14112 13499 14176
rect 13179 13088 13499 14112
rect 13179 13024 13187 13088
rect 13251 13024 13267 13088
rect 13331 13024 13347 13088
rect 13411 13024 13427 13088
rect 13491 13024 13499 13088
rect 13179 12000 13499 13024
rect 13179 11936 13187 12000
rect 13251 11936 13267 12000
rect 13331 11936 13347 12000
rect 13411 11936 13427 12000
rect 13491 11936 13499 12000
rect 13179 10912 13499 11936
rect 13179 10848 13187 10912
rect 13251 10848 13267 10912
rect 13331 10848 13347 10912
rect 13411 10848 13427 10912
rect 13491 10848 13499 10912
rect 13179 9824 13499 10848
rect 13179 9760 13187 9824
rect 13251 9760 13267 9824
rect 13331 9760 13347 9824
rect 13411 9760 13427 9824
rect 13491 9760 13499 9824
rect 13179 8736 13499 9760
rect 13179 8672 13187 8736
rect 13251 8672 13267 8736
rect 13331 8672 13347 8736
rect 13411 8672 13427 8736
rect 13491 8672 13499 8736
rect 13179 7648 13499 8672
rect 13179 7584 13187 7648
rect 13251 7584 13267 7648
rect 13331 7584 13347 7648
rect 13411 7584 13427 7648
rect 13491 7584 13499 7648
rect 13179 6560 13499 7584
rect 13179 6496 13187 6560
rect 13251 6496 13267 6560
rect 13331 6496 13347 6560
rect 13411 6496 13427 6560
rect 13491 6496 13499 6560
rect 13179 5472 13499 6496
rect 13179 5408 13187 5472
rect 13251 5408 13267 5472
rect 13331 5408 13347 5472
rect 13411 5408 13427 5472
rect 13491 5408 13499 5472
rect 13179 4384 13499 5408
rect 13179 4320 13187 4384
rect 13251 4320 13267 4384
rect 13331 4320 13347 4384
rect 13411 4320 13427 4384
rect 13491 4320 13499 4384
rect 13179 3296 13499 4320
rect 13179 3232 13187 3296
rect 13251 3232 13267 3296
rect 13331 3232 13347 3296
rect 13411 3232 13427 3296
rect 13491 3232 13499 3296
rect 13179 2208 13499 3232
rect 13179 2144 13187 2208
rect 13251 2144 13267 2208
rect 13331 2144 13347 2208
rect 13411 2144 13427 2208
rect 13491 2144 13499 2208
rect 13179 2128 13499 2144
use sky130_fd_sc_hd__inv_2  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 12144 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1717180972
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1717180972
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1717180972
transform -1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1717180972
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9844 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _167_
timestamp 1717180972
transform 1 0 10396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _168_
timestamp 1717180972
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1717180972
transform -1 0 12696 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _172_
timestamp 1717180972
transform -1 0 12052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1717180972
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _176_
timestamp 1717180972
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9568 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 8556 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 7452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6624 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _183_
timestamp 1717180972
transform 1 0 7268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _184_
timestamp 1717180972
transform 1 0 7820 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp 1717180972
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _187_
timestamp 1717180972
transform 1 0 6992 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _188_
timestamp 1717180972
transform 1 0 7176 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1717180972
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1717180972
transform -1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6808 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1717180972
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1717180972
transform 1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _194_
timestamp 1717180972
transform 1 0 5888 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _195_
timestamp 1717180972
transform -1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1717180972
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _197_
timestamp 1717180972
transform -1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6440 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _200_
timestamp 1717180972
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _201_
timestamp 1717180972
transform 1 0 6716 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 10488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp 1717180972
transform -1 0 3496 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _205_
timestamp 1717180972
transform -1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _206_
timestamp 1717180972
transform 1 0 9292 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1717180972
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1717180972
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _210_
timestamp 1717180972
transform 1 0 10488 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1717180972
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1717180972
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _213_
timestamp 1717180972
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _214_
timestamp 1717180972
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _215_
timestamp 1717180972
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _216_
timestamp 1717180972
transform -1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3404 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1717180972
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _219_
timestamp 1717180972
transform 1 0 3680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _220_
timestamp 1717180972
transform -1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3680 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1717180972
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _223_
timestamp 1717180972
transform -1 0 6164 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1717180972
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7360 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1717180972
transform -1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1717180972
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _229_
timestamp 1717180972
transform 1 0 8188 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9752 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1717180972
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _233_
timestamp 1717180972
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _234_
timestamp 1717180972
transform 1 0 9568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 1717180972
transform -1 0 11224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1717180972
transform 1 0 10948 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1717180972
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _239_
timestamp 1717180972
transform -1 0 10212 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 1717180972
transform 1 0 9936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _241_
timestamp 1717180972
transform 1 0 10212 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1717180972
transform -1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _243_
timestamp 1717180972
transform 1 0 7544 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _244_
timestamp 1717180972
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp 1717180972
transform -1 0 9752 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1717180972
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _247_
timestamp 1717180972
transform 1 0 8188 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _248_
timestamp 1717180972
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1717180972
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1717180972
transform -1 0 4324 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _251_
timestamp 1717180972
transform 1 0 5060 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _252_
timestamp 1717180972
transform 1 0 5336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1717180972
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _254_
timestamp 1717180972
transform 1 0 3312 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _255_
timestamp 1717180972
transform 1 0 4140 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _256_
timestamp 1717180972
transform 1 0 3956 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1717180972
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _258_
timestamp 1717180972
transform -1 0 4232 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _259_
timestamp 1717180972
transform -1 0 3404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1717180972
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _261_
timestamp 1717180972
transform -1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _263_
timestamp 1717180972
transform -1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1717180972
transform 1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1717180972
transform -1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1717180972
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _267_
timestamp 1717180972
transform -1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1717180972
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _269_
timestamp 1717180972
transform -1 0 2576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9016 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _271_
timestamp 1717180972
transform 1 0 9844 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _272_
timestamp 1717180972
transform 1 0 9108 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _274_
timestamp 1717180972
transform 1 0 9752 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _275_
timestamp 1717180972
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _276_
timestamp 1717180972
transform -1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _277_
timestamp 1717180972
transform 1 0 1932 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _278_
timestamp 1717180972
transform 1 0 2852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _279_
timestamp 1717180972
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _280_
timestamp 1717180972
transform -1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp 1717180972
transform 1 0 5060 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _282_
timestamp 1717180972
transform 1 0 5888 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _283_
timestamp 1717180972
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _285_
timestamp 1717180972
transform -1 0 8832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1717180972
transform -1 0 8004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _287_
timestamp 1717180972
transform 1 0 8924 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 1717180972
transform 1 0 8004 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _289_
timestamp 1717180972
transform 1 0 10672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 8832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _291_
timestamp 1717180972
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1717180972
transform -1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1717180972
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1717180972
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1717180972
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1717180972
transform -1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1717180972
transform -1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1717180972
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1717180972
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1717180972
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1717180972
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _303_
timestamp 1717180972
transform 1 0 2668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1717180972
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1717180972
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1717180972
transform 1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1717180972
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1717180972
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1717180972
transform 1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1717180972
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1717180972
transform 1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1717180972
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1717180972
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5428 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1717180972
transform -1 0 8280 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1717180972
transform 1 0 7728 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1717180972
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _319_
timestamp 1717180972
transform 1 0 2576 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _320_
timestamp 1717180972
transform 1 0 1472 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _321_
timestamp 1717180972
transform 1 0 4324 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1717180972
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _323_
timestamp 1717180972
transform -1 0 9108 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1717180972
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1717180972
transform 1 0 11132 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1717180972
transform 1 0 11132 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1717180972
transform 1 0 11132 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _328_
timestamp 1717180972
transform 1 0 5060 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3772 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _330_
timestamp 1717180972
transform 1 0 5060 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 1717180972
transform 1 0 7452 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _332_
timestamp 1717180972
transform 1 0 10212 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1717180972
transform 1 0 11132 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1717180972
transform -1 0 6440 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1717180972
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19
timestamp 1717180972
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 4416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_48
timestamp 1717180972
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57
timestamp 1717180972
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_63
timestamp 1717180972
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_70
timestamp 1717180972
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1717180972
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_88
timestamp 1717180972
transform 1 0 9200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1717180972
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104
timestamp 1717180972
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_123
timestamp 1717180972
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1717180972
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1717180972
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_42
timestamp 1717180972
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1717180972
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1717180972
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_64
timestamp 1717180972
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_75
timestamp 1717180972
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_84
timestamp 1717180972
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_94
timestamp 1717180972
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_113
timestamp 1717180972
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_119
timestamp 1717180972
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_126
timestamp 1717180972
transform 1 0 12696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_38
timestamp 1717180972
transform 1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_59
timestamp 1717180972
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_100
timestamp 1717180972
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_104
timestamp 1717180972
transform 1 0 10672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_129
timestamp 1717180972
transform 1 0 12972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1717180972
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1717180972
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_18
timestamp 1717180972
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_25
timestamp 1717180972
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_34
timestamp 1717180972
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1717180972
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1717180972
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_91
timestamp 1717180972
transform 1 0 9476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_97
timestamp 1717180972
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1717180972
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_120
timestamp 1717180972
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_6
timestamp 1717180972
transform 1 0 1656 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_14
timestamp 1717180972
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 1717180972
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1717180972
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1717180972
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1717180972
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1717180972
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1717180972
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1717180972
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1717180972
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1717180972
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 1717180972
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_103
timestamp 1717180972
transform 1 0 10580 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_107
timestamp 1717180972
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_129
timestamp 1717180972
transform 1 0 12972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1717180972
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_17
timestamp 1717180972
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_25
timestamp 1717180972
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_34
timestamp 1717180972
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1717180972
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1717180972
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_65
timestamp 1717180972
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_84
timestamp 1717180972
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_90
timestamp 1717180972
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_95
timestamp 1717180972
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_116
timestamp 1717180972
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_123
timestamp 1717180972
transform 1 0 12420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_129
timestamp 1717180972
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1717180972
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1717180972
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1717180972
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1717180972
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1717180972
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1717180972
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1717180972
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_121
timestamp 1717180972
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_129
timestamp 1717180972
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1717180972
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_11
timestamp 1717180972
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_20
timestamp 1717180972
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_29
timestamp 1717180972
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1717180972
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1717180972
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_82
timestamp 1717180972
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_88
timestamp 1717180972
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_101
timestamp 1717180972
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1717180972
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1717180972
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1717180972
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1717180972
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1717180972
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_38
timestamp 1717180972
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_42
timestamp 1717180972
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_68
timestamp 1717180972
transform 1 0 7360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1717180972
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1717180972
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_129
timestamp 1717180972
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1717180972
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1717180972
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 1717180972
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 1717180972
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_43
timestamp 1717180972
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1717180972
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_62
timestamp 1717180972
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 1717180972
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1717180972
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 1717180972
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1717180972
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_123
timestamp 1717180972
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_129
timestamp 1717180972
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1717180972
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_11
timestamp 1717180972
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1717180972
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1717180972
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 1717180972
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 1717180972
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1717180972
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1717180972
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_90
timestamp 1717180972
transform 1 0 9384 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_94
timestamp 1717180972
transform 1 0 9752 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_106
timestamp 1717180972
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_129
timestamp 1717180972
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1717180972
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1717180972
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_37
timestamp 1717180972
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_49
timestamp 1717180972
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_77
timestamp 1717180972
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_89
timestamp 1717180972
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1717180972
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1717180972
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_113
timestamp 1717180972
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1717180972
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 1717180972
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_46
timestamp 1717180972
transform 1 0 5336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_75
timestamp 1717180972
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1717180972
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1717180972
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1717180972
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_109
timestamp 1717180972
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_114
timestamp 1717180972
transform 1 0 11592 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_123
timestamp 1717180972
transform 1 0 12420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_129
timestamp 1717180972
transform 1 0 12972 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1717180972
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1717180972
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1717180972
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1717180972
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1717180972
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1717180972
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_70
timestamp 1717180972
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_92
timestamp 1717180972
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_97
timestamp 1717180972
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_101
timestamp 1717180972
transform 1 0 10396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1717180972
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_120
timestamp 1717180972
transform 1 0 12144 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_128
timestamp 1717180972
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1717180972
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_15
timestamp 1717180972
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_21
timestamp 1717180972
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1717180972
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1717180972
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_41
timestamp 1717180972
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_69
timestamp 1717180972
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1717180972
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1717180972
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_107
timestamp 1717180972
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_111
timestamp 1717180972
transform 1 0 11316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_126
timestamp 1717180972
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1717180972
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1717180972
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1717180972
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_35
timestamp 1717180972
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_41
timestamp 1717180972
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_49
timestamp 1717180972
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_63
timestamp 1717180972
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_81
timestamp 1717180972
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_89
timestamp 1717180972
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_102
timestamp 1717180972
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1717180972
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1717180972
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1717180972
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_59
timestamp 1717180972
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_69
timestamp 1717180972
transform 1 0 7452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_75
timestamp 1717180972
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1717180972
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1717180972
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_93
timestamp 1717180972
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_105
timestamp 1717180972
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_111
timestamp 1717180972
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_123
timestamp 1717180972
transform 1 0 12420 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_129
timestamp 1717180972
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1717180972
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1717180972
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1717180972
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_35
timestamp 1717180972
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_41
timestamp 1717180972
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1717180972
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 1717180972
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_68
timestamp 1717180972
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_80
timestamp 1717180972
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_102
timestamp 1717180972
transform 1 0 10488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_123
timestamp 1717180972
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_129
timestamp 1717180972
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1717180972
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1717180972
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1717180972
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1717180972
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 1717180972
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_64
timestamp 1717180972
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_71
timestamp 1717180972
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1717180972
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1717180972
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_101
timestamp 1717180972
transform 1 0 10396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_119
timestamp 1717180972
transform 1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_127
timestamp 1717180972
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1717180972
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1717180972
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1717180972
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1717180972
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1717180972
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1717180972
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_62
timestamp 1717180972
transform 1 0 6808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_90
timestamp 1717180972
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_97
timestamp 1717180972
transform 1 0 10028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_101
timestamp 1717180972
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1717180972
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1717180972
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_116
timestamp 1717180972
transform 1 0 11776 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1717180972
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1717180972
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1717180972
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1717180972
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1717180972
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1717180972
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1717180972
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_65
timestamp 1717180972
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_70
timestamp 1717180972
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1717180972
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1717180972
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_90
timestamp 1717180972
transform 1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_96
timestamp 1717180972
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_120
timestamp 1717180972
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_128
timestamp 1717180972
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1717180972
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1717180972
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_27
timestamp 1717180972
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_35
timestamp 1717180972
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1717180972
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1717180972
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1717180972
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1717180972
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_81
timestamp 1717180972
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_85
timestamp 1717180972
transform 1 0 8924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_97
timestamp 1717180972
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_105
timestamp 1717180972
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1717180972
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_125
timestamp 1717180972
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1717180972
transform -1 0 13064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1717180972
transform 1 0 7360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1717180972
transform -1 0 13064 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1717180972
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1717180972
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1717180972
transform 1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1717180972
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1717180972
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1717180972
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1717180972
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1717180972
transform -1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1717180972
transform -1 0 13064 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1717180972
transform -1 0 13064 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1717180972
transform -1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1717180972
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 4324 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1717180972
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1717180972
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1717180972
transform -1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1717180972
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1717180972
transform -1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1717180972
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1717180972
transform -1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1717180972
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1717180972
transform -1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1717180972
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1717180972
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1717180972
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1717180972
transform -1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1717180972
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1717180972
transform -1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1717180972
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1717180972
transform -1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1717180972
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1717180972
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1717180972
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1717180972
transform -1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1717180972
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1717180972
transform -1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1717180972
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1717180972
transform -1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1717180972
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1717180972
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1717180972
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1717180972
transform -1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1717180972
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1717180972
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1717180972
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1717180972
transform -1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1717180972
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1717180972
transform -1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1717180972
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1717180972
transform -1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1717180972
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1717180972
transform -1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1717180972
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1717180972
transform -1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1717180972
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1717180972
transform -1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1717180972
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1717180972
transform -1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1717180972
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1717180972
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1717180972
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1717180972
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1717180972
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1717180972
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1717180972
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1717180972
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1717180972
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1717180972
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1717180972
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1717180972
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1717180972
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1717180972
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1717180972
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1717180972
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1717180972
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1717180972
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1717180972
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1717180972
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1717180972
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1717180972
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1717180972
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1717180972
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1717180972
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1717180972
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1717180972
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1717180972
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1717180972
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1717180972
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1717180972
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1717180972
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1717180972
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1717180972
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1717180972
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1717180972
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1717180972
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1717180972
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1717180972
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1717180972
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1717180972
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1717180972
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1717180972
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1717180972
transform 1 0 3680 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1717180972
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1717180972
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1717180972
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 4002 2128 4322 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7061 2128 7381 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10120 2128 10440 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 13179 2128 13499 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2473 2128 2793 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5532 2128 5852 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8591 2128 8911 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11650 2128 11970 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 pulse_count[0]
port 3 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 pulse_count[1]
port 4 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 pulse_count[2]
port 5 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 pulse_count[3]
port 6 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 pulse_count[4]
port 7 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 pulse_count[5]
port 8 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 pulse_count[6]
port 9 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 pulse_count[7]
port 10 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 pulse_count[8]
port 11 nsew signal input
flabel metal3 s 13657 1912 14457 2032 0 FreeSans 480 0 0 0 pulse_period[0]
port 12 nsew signal input
flabel metal3 s 13657 5992 14457 6112 0 FreeSans 480 0 0 0 pulse_period[1]
port 13 nsew signal input
flabel metal3 s 13657 10072 14457 10192 0 FreeSans 480 0 0 0 pulse_period[2]
port 14 nsew signal input
flabel metal3 s 13657 14152 14457 14272 0 FreeSans 480 0 0 0 pulse_period[3]
port 15 nsew signal input
flabel metal2 s 3606 15801 3662 16601 0 FreeSans 224 90 0 0 pwm_out1
port 16 nsew signal tristate
flabel metal2 s 10782 15801 10838 16601 0 FreeSans 224 90 0 0 pwm_out2
port 17 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 rst
port 18 nsew signal input
rlabel via1 7301 14144 7301 14144 0 VGND
rlabel metal1 7222 13600 7222 13600 0 VPWR
rlabel metal1 7137 8942 7137 8942 0 _000_
rlabel metal1 7551 5610 7551 5610 0 _001_
rlabel metal1 8418 9146 8418 9146 0 _002_
rlabel metal1 3135 6698 3135 6698 0 _003_
rlabel metal1 2583 8874 2583 8874 0 _004_
rlabel metal1 4377 9622 4377 9622 0 _005_
rlabel metal2 2898 5882 2898 5882 0 _006_
rlabel metal1 5842 5338 5842 5338 0 _007_
rlabel metal1 6624 7174 6624 7174 0 _008_
rlabel metal2 8050 7582 8050 7582 0 _009_
rlabel metal1 10955 7446 10955 7446 0 _010_
rlabel metal1 12236 7174 12236 7174 0 _011_
rlabel metal2 12190 4760 12190 4760 0 _012_
rlabel metal2 12558 3332 12558 3332 0 _013_
rlabel metal2 6026 9826 6026 9826 0 _014_
rlabel metal2 4738 10914 4738 10914 0 _015_
rlabel metal1 5888 12682 5888 12682 0 _016_
rlabel metal1 8556 12410 8556 12410 0 _017_
rlabel metal2 11638 13124 11638 13124 0 _018_
rlabel metal2 12190 8024 12190 8024 0 _019_
rlabel metal2 5750 8738 5750 8738 0 _020_
rlabel metal1 8381 5882 8381 5882 0 _021_
rlabel metal1 8050 9656 8050 9656 0 _022_
rlabel metal1 1971 6970 1971 6970 0 _023_
rlabel metal1 3128 8602 3128 8602 0 _024_
rlabel metal1 3036 9622 3036 9622 0 _025_
rlabel metal1 1978 5746 1978 5746 0 _026_
rlabel metal1 4692 6358 4692 6358 0 _027_
rlabel metal1 5888 6834 5888 6834 0 _028_
rlabel metal1 8602 7446 8602 7446 0 _029_
rlabel metal2 9522 7582 9522 7582 0 _030_
rlabel metal1 11270 6698 11270 6698 0 _031_
rlabel metal1 11500 4658 11500 4658 0 _032_
rlabel metal1 12236 3162 12236 3162 0 _033_
rlabel metal2 5934 10268 5934 10268 0 _034_
rlabel metal1 4363 11322 4363 11322 0 _035_
rlabel via1 5658 12155 5658 12155 0 _036_
rlabel metal1 7820 12886 7820 12886 0 _037_
rlabel metal1 10212 13226 10212 13226 0 _038_
rlabel metal2 11454 8364 11454 8364 0 _039_
rlabel metal1 6992 12886 6992 12886 0 _040_
rlabel metal1 7452 12410 7452 12410 0 _041_
rlabel metal1 8786 12342 8786 12342 0 _042_
rlabel metal1 9522 13294 9522 13294 0 _043_
rlabel metal1 7368 12138 7368 12138 0 _044_
rlabel metal1 7866 12410 7866 12410 0 _045_
rlabel metal1 6900 11866 6900 11866 0 _046_
rlabel metal1 6762 11322 6762 11322 0 _047_
rlabel metal1 6256 12818 6256 12818 0 _048_
rlabel metal1 6762 10710 6762 10710 0 _049_
rlabel metal1 6164 10778 6164 10778 0 _050_
rlabel metal1 7590 10506 7590 10506 0 _051_
rlabel metal2 6946 3298 6946 3298 0 _052_
rlabel metal1 7268 3706 7268 3706 0 _053_
rlabel metal1 10471 4114 10471 4114 0 _054_
rlabel metal1 5106 9078 5106 9078 0 _055_
rlabel metal1 2346 8398 2346 8398 0 _056_
rlabel metal1 4692 5270 4692 5270 0 _057_
rlabel metal1 5198 7242 5198 7242 0 _058_
rlabel metal1 10074 5202 10074 5202 0 _059_
rlabel metal1 11132 5270 11132 5270 0 _060_
rlabel metal1 12144 3026 12144 3026 0 _061_
rlabel metal1 11040 4998 11040 4998 0 _062_
rlabel metal1 9890 3502 9890 3502 0 _063_
rlabel metal1 5198 3536 5198 3536 0 _064_
rlabel metal1 4186 3638 4186 3638 0 _065_
rlabel metal1 2944 3162 2944 3162 0 _066_
rlabel metal1 1886 3400 1886 3400 0 _067_
rlabel metal2 3082 3332 3082 3332 0 _068_
rlabel metal1 5014 3536 5014 3536 0 _069_
rlabel metal1 4094 3604 4094 3604 0 _070_
rlabel metal1 4278 3060 4278 3060 0 _071_
rlabel metal1 4554 3026 4554 3026 0 _072_
rlabel metal1 4416 2822 4416 2822 0 _073_
rlabel metal1 6486 2414 6486 2414 0 _074_
rlabel metal1 5658 3094 5658 3094 0 _075_
rlabel metal1 6210 3706 6210 3706 0 _076_
rlabel metal1 7728 3366 7728 3366 0 _077_
rlabel metal1 8878 4046 8878 4046 0 _078_
rlabel metal1 8786 3570 8786 3570 0 _079_
rlabel metal1 9476 3502 9476 3502 0 _080_
rlabel metal1 8970 3162 8970 3162 0 _081_
rlabel metal1 9430 3434 9430 3434 0 _082_
rlabel metal2 9706 3332 9706 3332 0 _083_
rlabel metal1 10948 3706 10948 3706 0 _084_
rlabel metal1 9614 3536 9614 3536 0 _085_
rlabel metal1 10488 3706 10488 3706 0 _086_
rlabel metal1 10810 4012 10810 4012 0 _087_
rlabel metal1 2254 7956 2254 7956 0 _088_
rlabel metal1 11546 5202 11546 5202 0 _089_
rlabel metal1 9890 6358 9890 6358 0 _090_
rlabel metal1 10488 6426 10488 6426 0 _091_
rlabel metal1 10856 6766 10856 6766 0 _092_
rlabel metal1 8510 6766 8510 6766 0 _093_
rlabel metal2 9338 7208 9338 7208 0 _094_
rlabel metal1 9200 6970 9200 6970 0 _095_
rlabel metal1 8510 6426 8510 6426 0 _096_
rlabel metal1 8556 6970 8556 6970 0 _097_
rlabel metal1 4186 6426 4186 6426 0 _098_
rlabel metal2 6118 7072 6118 7072 0 _099_
rlabel metal1 6072 7378 6072 7378 0 _100_
rlabel metal1 3542 6086 3542 6086 0 _101_
rlabel metal1 4462 5610 4462 5610 0 _102_
rlabel metal1 4738 5882 4738 5882 0 _103_
rlabel metal1 3404 5270 3404 5270 0 _104_
rlabel metal1 2691 6290 2691 6290 0 _105_
rlabel metal1 2484 8466 2484 8466 0 _106_
rlabel metal1 3772 8534 3772 8534 0 _107_
rlabel metal2 3358 9316 3358 9316 0 _108_
rlabel metal1 2530 7888 2530 7888 0 _109_
rlabel metal1 2622 8500 2622 8500 0 _110_
rlabel metal1 2576 7514 2576 7514 0 _111_
rlabel metal1 9200 11322 9200 11322 0 _112_
rlabel metal1 9522 11866 9522 11866 0 _113_
rlabel metal1 9752 12410 9752 12410 0 _114_
rlabel metal1 10258 12240 10258 12240 0 _115_
rlabel metal1 9108 10642 9108 10642 0 _116_
rlabel metal1 4692 3162 4692 3162 0 _117_
rlabel metal1 3266 3536 3266 3536 0 _118_
rlabel metal1 3818 3536 3818 3536 0 _119_
rlabel metal1 4692 3706 4692 3706 0 _120_
rlabel metal1 5428 4114 5428 4114 0 _121_
rlabel metal1 5796 3162 5796 3162 0 _122_
rlabel metal1 5980 3570 5980 3570 0 _123_
rlabel metal1 7130 3094 7130 3094 0 _124_
rlabel metal2 7498 3196 7498 3196 0 _125_
rlabel metal1 7774 3060 7774 3060 0 _126_
rlabel metal1 8050 3162 8050 3162 0 _127_
rlabel metal1 8510 3706 8510 3706 0 _128_
rlabel metal1 8556 4250 8556 4250 0 _129_
rlabel metal1 9982 4794 9982 4794 0 _130_
rlabel metal1 2944 6290 2944 6290 0 _131_
rlabel metal2 5244 8398 5244 8398 0 _132_
rlabel metal1 12328 9146 12328 9146 0 _133_
rlabel metal1 7452 4250 7452 4250 0 _134_
rlabel metal1 10534 11526 10534 11526 0 _135_
rlabel metal2 9522 10948 9522 10948 0 _136_
rlabel metal1 10120 12682 10120 12682 0 _137_
rlabel metal1 10074 11696 10074 11696 0 _138_
rlabel via1 8313 5270 8313 5270 0 _139_
rlabel metal2 9798 10438 9798 10438 0 _140_
rlabel metal1 10166 9894 10166 9894 0 _141_
rlabel metal1 10764 10234 10764 10234 0 _142_
rlabel metal1 11454 10506 11454 10506 0 _143_
rlabel metal1 12098 10098 12098 10098 0 _144_
rlabel metal1 11960 10778 11960 10778 0 _145_
rlabel metal1 11960 10506 11960 10506 0 _146_
rlabel metal1 11454 11662 11454 11662 0 _147_
rlabel metal1 9982 10676 9982 10676 0 _148_
rlabel metal1 12006 11152 12006 11152 0 _149_
rlabel metal1 10764 9690 10764 9690 0 _150_
rlabel metal1 11362 10030 11362 10030 0 _151_
rlabel metal1 12144 10234 12144 10234 0 _152_
rlabel metal1 10074 10608 10074 10608 0 _153_
rlabel metal1 9016 10710 9016 10710 0 _154_
rlabel metal2 6762 13124 6762 13124 0 _155_
rlabel metal1 6624 10642 6624 10642 0 _156_
rlabel metal2 4094 12189 4094 12189 0 clk
rlabel metal1 7360 7854 7360 7854 0 clknet_0_clk
rlabel metal2 11178 4080 11178 4080 0 clknet_1_0__leaf_clk
rlabel metal1 2622 9418 2622 9418 0 clknet_1_1__leaf_clk
rlabel metal1 2346 3638 2346 3638 0 counter1\[0\]
rlabel metal1 12926 4148 12926 4148 0 counter1\[10\]
rlabel metal1 2208 3366 2208 3366 0 counter1\[1\]
rlabel metal1 4311 8942 4311 8942 0 counter1\[2\]
rlabel metal1 4554 4148 4554 4148 0 counter1\[3\]
rlabel metal1 4324 6358 4324 6358 0 counter1\[4\]
rlabel metal2 5566 5389 5566 5389 0 counter1\[5\]
rlabel metal2 7636 4114 7636 4114 0 counter1\[6\]
rlabel metal1 9430 5202 9430 5202 0 counter1\[7\]
rlabel metal1 9798 5270 9798 5270 0 counter1\[8\]
rlabel metal1 11178 4250 11178 4250 0 counter1\[9\]
rlabel metal1 9706 9588 9706 9588 0 counter2\[0\]
rlabel metal1 9384 11118 9384 11118 0 counter2\[1\]
rlabel metal1 11776 10574 11776 10574 0 counter2\[2\]
rlabel metal1 10074 12138 10074 12138 0 counter2\[3\]
rlabel metal1 10350 12274 10350 12274 0 counter2\[4\]
rlabel metal2 12926 8228 12926 8228 0 counter2\[5\]
rlabel metal1 2116 3638 2116 3638 0 net1
rlabel metal1 12788 2618 12788 2618 0 net10
rlabel metal1 12650 10234 12650 10234 0 net11
rlabel metal1 11500 9622 11500 9622 0 net12
rlabel metal1 10718 12852 10718 12852 0 net13
rlabel via1 2162 4590 2162 4590 0 net14
rlabel metal1 6394 5882 6394 5882 0 net15
rlabel metal1 10810 9520 10810 9520 0 net16
rlabel metal2 6118 8806 6118 8806 0 net17
rlabel metal2 12374 8772 12374 8772 0 net18
rlabel metal1 8096 5134 8096 5134 0 net19
rlabel metal1 3266 2618 3266 2618 0 net2
rlabel metal1 12052 4114 12052 4114 0 net20
rlabel metal1 7912 10642 7912 10642 0 net21
rlabel metal1 4646 2618 4646 2618 0 net3
rlabel metal1 6026 2618 6026 2618 0 net4
rlabel metal1 6486 2584 6486 2584 0 net5
rlabel metal1 8786 3026 8786 3026 0 net6
rlabel metal1 10074 2618 10074 2618 0 net7
rlabel metal1 8418 3468 8418 3468 0 net8
rlabel metal2 10902 3196 10902 3196 0 net9
rlabel metal1 5014 8942 5014 8942 0 prev_pwm_out2
rlabel metal2 966 1588 966 1588 0 pulse_count[0]
rlabel metal2 2530 1027 2530 1027 0 pulse_count[1]
rlabel metal2 4094 1027 4094 1027 0 pulse_count[2]
rlabel metal2 5658 1027 5658 1027 0 pulse_count[3]
rlabel metal2 7222 823 7222 823 0 pulse_count[4]
rlabel metal2 8786 1588 8786 1588 0 pulse_count[5]
rlabel metal2 10350 823 10350 823 0 pulse_count[6]
rlabel metal2 11914 1554 11914 1554 0 pulse_count[7]
rlabel metal2 13478 1163 13478 1163 0 pulse_count[8]
rlabel metal1 12972 2346 12972 2346 0 pulse_period[0]
rlabel metal2 13018 6137 13018 6137 0 pulse_period[1]
rlabel metal2 13018 10353 13018 10353 0 pulse_period[2]
rlabel metal1 13110 13974 13110 13974 0 pulse_period[3]
rlabel metal1 3772 14042 3772 14042 0 pwm_out1
rlabel metal2 10810 14936 10810 14936 0 pwm_out2
rlabel metal3 820 4148 820 4148 0 rst
<< properties >>
string FIXED_BBOX 0 0 14457 16601
<< end >>
