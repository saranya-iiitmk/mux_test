magic
tech sky130A
timestamp 1717060164
use sky130_fd_pr__cap_mim_m3_1_P9YBYH  XC2
timestamp 1717060164
transform 1 0 193 0 1 1820
box -193 -1520 193 1520
<< end >>
