magic
tech sky130A
magscale 1 2
timestamp 1717180972
<< nwell >>
rect -508 998 -330 1064
rect -138 1016 158 1064
rect -112 998 154 1016
rect -508 928 612 998
rect -508 729 508 928
rect 746 738 1067 1062
rect 1431 768 1432 860
rect 1736 754 1766 768
rect -508 719 511 729
rect -508 707 518 719
rect -508 699 533 707
rect -508 684 518 699
rect -508 658 252 684
rect -508 494 108 658
rect 488 624 518 684
rect 612 678 1067 738
rect 612 677 746 678
rect 740 620 774 657
rect -508 371 256 494
rect -110 362 256 371
rect -1 360 256 362
rect -1 355 12 360
rect 822 354 1067 678
rect 1678 739 1711 741
rect 1735 739 1766 754
rect 1870 739 1887 754
rect 1554 642 1584 672
rect 1678 666 2070 739
rect 1678 354 1711 666
rect 1805 630 1835 639
<< psubdiff >>
rect -890 882 -744 921
rect -890 788 -849 882
rect -780 788 -744 882
rect -890 738 -744 788
<< nsubdiff >>
rect -455 799 -351 823
rect -455 749 -429 799
rect -376 749 -351 799
rect -455 721 -351 749
<< psubdiffcont >>
rect -849 788 -780 882
<< nsubdiffcont >>
rect -429 749 -376 799
<< poly >>
rect -236 1632 366 1662
rect -236 1433 -206 1632
rect 36 1572 106 1589
rect 36 1537 52 1572
rect 89 1567 106 1572
rect 89 1537 278 1567
rect 36 1533 278 1537
rect 36 1517 106 1533
rect 248 1483 278 1533
rect 336 1492 366 1632
rect 1314 1618 1766 1648
rect 1314 1497 1344 1618
rect 1587 1532 1653 1548
rect 1587 1530 1603 1532
rect 1402 1500 1603 1530
rect 1402 1498 1432 1500
rect 1587 1498 1603 1500
rect 1637 1498 1653 1532
rect 1587 1482 1653 1498
rect 1736 1360 1766 1618
rect 1402 1098 1566 1128
rect 1536 1094 1566 1098
rect 1536 1064 1766 1094
rect 55 820 127 838
rect 55 785 75 820
rect 110 813 127 820
rect 336 813 366 865
rect 110 785 366 813
rect 55 776 366 785
rect 55 766 127 776
rect 1736 754 1900 784
rect -61 719 5 733
rect 1870 732 1900 754
rect -61 682 -45 719
rect -11 688 518 719
rect -11 682 5 688
rect -61 649 5 682
rect 182 640 212 688
rect 488 624 518 688
rect 1248 700 1584 730
rect 1248 637 1278 700
rect 1554 661 1584 700
rect 1870 722 1950 732
rect 1870 688 1900 722
rect 1934 688 1950 722
rect 1877 678 1950 688
rect 1554 631 1835 661
rect 1805 615 1835 631
rect 1666 346 1732 362
rect 1666 326 1682 346
rect 1278 296 1466 326
rect 1584 312 1682 326
rect 1716 312 1732 346
rect 1584 296 1732 312
rect -234 -361 -204 76
rect -107 -33 -40 -16
rect -107 -67 -94 -33
rect -55 -67 -40 -33
rect -107 -85 -40 -67
rect -83 -196 -53 -85
rect 94 -196 124 0
rect 182 -57 212 8
rect 182 -68 256 -57
rect 182 -102 205 -68
rect 240 -102 256 -68
rect 182 -138 256 -102
rect 400 -196 430 26
rect -83 -226 430 -196
rect 180 -357 262 -337
rect 180 -361 206 -357
rect -234 -391 206 -361
rect 241 -361 262 -357
rect 488 -361 518 12
rect 1160 -73 1190 2
rect 1466 -50 1496 1
rect 1805 -50 1835 44
rect 1953 -48 2019 -38
rect 1953 -50 1969 -48
rect 1466 -73 1969 -50
rect 1160 -80 1969 -73
rect 1160 -103 1496 -80
rect 1953 -82 1969 -80
rect 2003 -82 2019 -48
rect 1953 -92 2019 -82
rect 241 -391 518 -361
rect 180 -424 262 -391
<< polycont >>
rect 52 1537 89 1572
rect 1603 1498 1637 1532
rect 75 785 110 820
rect -45 682 -11 719
rect 1900 688 1934 722
rect 1682 312 1716 346
rect -94 -67 -55 -33
rect 205 -102 240 -68
rect 206 -391 241 -357
rect 1969 -82 2003 -48
<< locali >>
rect 36 1572 106 1589
rect 36 1567 52 1572
rect -194 1537 52 1567
rect 89 1537 106 1572
rect -194 1533 106 1537
rect -194 1417 -160 1533
rect 36 1517 106 1533
rect 290 1517 698 1551
rect -849 1274 -322 1308
rect -849 1272 -487 1274
rect -849 921 -775 1272
rect 290 1229 324 1517
rect 664 1337 698 1517
rect 1019 1549 1390 1583
rect -433 934 -328 970
rect -890 882 -744 921
rect -890 788 -849 882
rect -780 788 -744 882
rect -433 823 -394 934
rect -890 738 -744 788
rect -455 799 -351 823
rect -455 749 -429 799
rect -376 749 -351 799
rect -194 813 -160 880
rect 55 820 127 838
rect 55 813 75 820
rect -194 785 75 813
rect 110 785 127 820
rect -194 777 127 785
rect 55 766 127 777
rect -846 232 -776 738
rect -455 721 -351 749
rect -61 722 5 733
rect -432 573 -395 721
rect -192 719 5 722
rect -192 686 -45 719
rect -192 612 -158 686
rect -61 682 -45 686
rect -11 682 5 719
rect -61 649 5 682
rect 575 716 611 803
rect 575 680 775 716
rect 740 620 774 680
rect -432 536 -279 573
rect 1019 373 1053 1549
rect 1356 1475 1390 1549
rect 1587 1532 1653 1548
rect 1587 1498 1603 1532
rect 1637 1531 1653 1532
rect 1637 1498 1812 1531
rect 1587 1497 1812 1498
rect 1587 1482 1653 1497
rect 1778 1338 1812 1497
rect 1900 722 1934 1089
rect 1900 672 1934 688
rect 652 339 1053 373
rect 1666 346 1732 362
rect 1666 312 1682 346
rect 1716 312 1881 346
rect 1666 296 1732 312
rect -846 222 -308 232
rect -845 198 -308 222
rect -192 -34 -157 94
rect -107 -33 -40 -16
rect -107 -34 -94 -33
rect -192 -67 -94 -34
rect -55 -67 -40 -33
rect 1969 -48 2003 66
rect -192 -69 -40 -67
rect -107 -85 -40 -69
rect 182 -68 256 -57
rect 182 -102 205 -68
rect 240 -102 256 -68
rect 1969 -98 2003 -82
rect 182 -138 256 -102
rect 200 -337 235 -138
rect 180 -357 262 -337
rect 180 -391 206 -357
rect 241 -391 262 -357
rect 180 -424 262 -391
use inverter  inverter_0
timestamp 1717180972
transform 1 0 -280 0 1 -580
box -78 644 170 1266
use inverter  inverter_1
timestamp 1717180972
transform -1 0 698 0 -1 2004
box -78 644 170 1266
use inverter  inverter_2
timestamp 1717180972
transform 1 0 -282 0 -1 2086
box -78 644 170 1266
use inverter  inverter_3
timestamp 1717180972
transform -1 0 774 0 1 -588
box -78 644 170 1266
use inverter  inverter_4
timestamp 1717180972
transform -1 0 2022 0 -1 2004
box -78 644 170 1266
use inverter  inverter_5
timestamp 1717180972
transform 1 0 1690 0 -1 2004
box -78 644 170 1266
use inverter  inverter_6
timestamp 1717180972
transform 1 0 1759 0 1 -600
box -78 644 170 1266
use inverter  inverter_7
timestamp 1717180972
transform -1 0 2091 0 1 -600
box -78 644 170 1266
use mux1_4  mux1_4_0
timestamp 1717180972
transform 1 0 0 0 1 0
box 0 0 612 1498
use mux1_4  mux1_4_1
timestamp 1717180972
transform 1 0 1066 0 1 0
box 0 0 612 1498
<< end >>
