magic
tech sky130A
magscale 1 2
timestamp 1717237536
<< viali >>
rect 3249 11305 3283 11339
rect 9229 11305 9263 11339
rect 4629 11101 4663 11135
rect 3157 11033 3191 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 9137 11033 9171 11067
rect 4077 10965 4111 10999
rect 7297 10965 7331 10999
rect 2329 10761 2363 10795
rect 9045 10761 9079 10795
rect 5396 10693 5430 10727
rect 5733 10693 5767 10727
rect 1409 10625 1443 10659
rect 3065 10625 3099 10659
rect 3433 10625 3467 10659
rect 3617 10625 3651 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 8309 10625 8343 10659
rect 10425 10625 10459 10659
rect 3341 10557 3375 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 7021 10557 7055 10591
rect 8033 10557 8067 10591
rect 7113 10489 7147 10523
rect 1593 10421 1627 10455
rect 3525 10421 3559 10455
rect 4261 10421 4295 10455
rect 6377 10421 6411 10455
rect 10241 10421 10275 10455
rect 3249 10217 3283 10251
rect 3617 10217 3651 10251
rect 6101 10217 6135 10251
rect 7665 10217 7699 10251
rect 8401 10217 8435 10251
rect 9413 10217 9447 10251
rect 8125 10149 8159 10183
rect 3341 10081 3375 10115
rect 6285 10081 6319 10115
rect 8033 10081 8067 10115
rect 9597 10081 9631 10115
rect 2973 10013 3007 10047
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 9873 10013 9907 10047
rect 4046 9945 4080 9979
rect 6552 9945 6586 9979
rect 5181 9877 5215 9911
rect 5273 9877 5307 9911
rect 7757 9877 7791 9911
rect 9689 9877 9723 9911
rect 6561 9673 6595 9707
rect 6745 9673 6779 9707
rect 7665 9673 7699 9707
rect 8401 9673 8435 9707
rect 9312 9605 9346 9639
rect 3893 9537 3927 9571
rect 4169 9537 4203 9571
rect 5641 9537 5675 9571
rect 6742 9537 6776 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 8309 9537 8343 9571
rect 8585 9537 8619 9571
rect 4813 9469 4847 9503
rect 5089 9469 5123 9503
rect 7113 9469 7147 9503
rect 7205 9469 7239 9503
rect 9045 9469 9079 9503
rect 3617 9333 3651 9367
rect 4077 9333 4111 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 8125 9333 8159 9367
rect 10425 9333 10459 9367
rect 4905 9129 4939 9163
rect 5549 9129 5583 9163
rect 4261 8993 4295 9027
rect 10425 8993 10459 9027
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 9689 8925 9723 8959
rect 9781 8925 9815 8959
rect 6377 8857 6411 8891
rect 7665 8857 7699 8891
rect 7849 8857 7883 8891
rect 8033 8857 8067 8891
rect 5825 8789 5859 8823
rect 9597 8789 9631 8823
rect 7481 8585 7515 8619
rect 6561 8517 6595 8551
rect 6745 8517 6779 8551
rect 1593 8449 1627 8483
rect 4077 8449 4111 8483
rect 7297 8449 7331 8483
rect 7573 8449 7607 8483
rect 8197 8449 8231 8483
rect 1869 8381 1903 8415
rect 7941 8381 7975 8415
rect 3341 8313 3375 8347
rect 7113 8313 7147 8347
rect 3893 8245 3927 8279
rect 6377 8245 6411 8279
rect 9321 8245 9355 8279
rect 1593 8041 1627 8075
rect 7113 8041 7147 8075
rect 9873 8041 9907 8075
rect 2053 7905 2087 7939
rect 3065 7905 3099 7939
rect 3525 7905 3559 7939
rect 9505 7905 9539 7939
rect 1961 7837 1995 7871
rect 3433 7837 3467 7871
rect 7757 7837 7791 7871
rect 8585 7837 8619 7871
rect 9321 7837 9355 7871
rect 9781 7837 9815 7871
rect 9965 7837 9999 7871
rect 10057 7837 10091 7871
rect 10241 7837 10275 7871
rect 5273 7769 5307 7803
rect 6561 7701 6595 7735
rect 7941 7701 7975 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 10149 7701 10183 7735
rect 7757 7497 7791 7531
rect 8677 7497 8711 7531
rect 9505 7497 9539 7531
rect 8309 7429 8343 7463
rect 10333 7429 10367 7463
rect 1685 7361 1719 7395
rect 3801 7361 3835 7395
rect 5917 7361 5951 7395
rect 6377 7361 6411 7395
rect 6633 7361 6667 7395
rect 8769 7361 8803 7395
rect 8953 7361 8987 7395
rect 9413 7361 9447 7395
rect 10149 7361 10183 7395
rect 1961 7293 1995 7327
rect 4077 7293 4111 7327
rect 6193 7293 6227 7327
rect 8033 7293 8067 7327
rect 8217 7293 8251 7327
rect 9229 7293 9263 7327
rect 5733 7225 5767 7259
rect 3433 7157 3467 7191
rect 5549 7157 5583 7191
rect 6101 7157 6135 7191
rect 8953 7157 8987 7191
rect 9873 7157 9907 7191
rect 9965 7157 9999 7191
rect 1961 6953 1995 6987
rect 3985 6953 4019 6987
rect 8953 6953 8987 6987
rect 8769 6885 8803 6919
rect 2145 6817 2179 6851
rect 4997 6817 5031 6851
rect 5273 6817 5307 6851
rect 9505 6817 9539 6851
rect 10241 6817 10275 6851
rect 2237 6749 2271 6783
rect 3801 6749 3835 6783
rect 7389 6749 7423 6783
rect 5365 6681 5399 6715
rect 7656 6681 7690 6715
rect 6653 6613 6687 6647
rect 9689 6613 9723 6647
rect 7757 6409 7791 6443
rect 8953 6409 8987 6443
rect 10425 6409 10459 6443
rect 9290 6341 9324 6375
rect 3985 6273 4019 6307
rect 4629 6273 4663 6307
rect 6377 6273 6411 6307
rect 7941 6273 7975 6307
rect 8585 6273 8619 6307
rect 3893 6205 3927 6239
rect 4537 6205 4571 6239
rect 5089 6205 5123 6239
rect 8493 6205 8527 6239
rect 9045 6205 9079 6239
rect 4353 6137 4387 6171
rect 4997 6069 5031 6103
rect 5733 6069 5767 6103
rect 6561 6069 6595 6103
rect 1869 5865 1903 5899
rect 7297 5865 7331 5899
rect 8401 5865 8435 5899
rect 10057 5865 10091 5899
rect 2421 5797 2455 5831
rect 2237 5729 2271 5763
rect 2881 5729 2915 5763
rect 3341 5729 3375 5763
rect 3617 5729 3651 5763
rect 4077 5729 4111 5763
rect 5825 5729 5859 5763
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 3249 5661 3283 5695
rect 5457 5661 5491 5695
rect 5549 5661 5583 5695
rect 8677 5661 8711 5695
rect 9781 5661 9815 5695
rect 9965 5661 9999 5695
rect 10149 5661 10183 5695
rect 4721 5525 4755 5559
rect 5273 5525 5307 5559
rect 8217 5525 8251 5559
rect 9229 5525 9263 5559
rect 3985 5321 4019 5355
rect 5457 5253 5491 5287
rect 6653 5253 6687 5287
rect 8760 5253 8794 5287
rect 8493 5185 8527 5219
rect 1961 5117 1995 5151
rect 2237 5117 2271 5151
rect 5733 5117 5767 5151
rect 6377 5117 6411 5151
rect 3709 4981 3743 5015
rect 8125 4981 8159 5015
rect 9873 4981 9907 5015
rect 9321 4777 9355 4811
rect 9689 4777 9723 4811
rect 9229 4709 9263 4743
rect 4169 4641 4203 4675
rect 8677 4641 8711 4675
rect 9137 4641 9171 4675
rect 10333 4641 10367 4675
rect 4445 4573 4479 4607
rect 7297 4573 7331 4607
rect 8953 4573 8987 4607
rect 9413 4573 9447 4607
rect 9781 4573 9815 4607
rect 7941 4437 7975 4471
rect 8033 4437 8067 4471
rect 7205 4233 7239 4267
rect 8125 4233 8159 4267
rect 3341 4097 3375 4131
rect 4169 4097 4203 4131
rect 4629 4097 4663 4131
rect 7481 4097 7515 4131
rect 7573 4097 7607 4131
rect 7665 4097 7699 4131
rect 7941 4097 7975 4131
rect 8769 4097 8803 4131
rect 9781 4097 9815 4131
rect 3433 4029 3467 4063
rect 3709 4029 3743 4063
rect 4077 4029 4111 4063
rect 4537 4029 4571 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 8907 4029 8941 4063
rect 9045 4029 9079 4063
rect 9965 4029 9999 4063
rect 7757 3961 7791 3995
rect 9321 3961 9355 3995
rect 3801 3893 3835 3927
rect 5825 3893 5859 3927
rect 4537 3689 4571 3723
rect 5536 3689 5570 3723
rect 7021 3689 7055 3723
rect 8493 3689 8527 3723
rect 10425 3689 10459 3723
rect 1593 3553 1627 3587
rect 5273 3553 5307 3587
rect 7113 3553 7147 3587
rect 9045 3553 9079 3587
rect 4353 3485 4387 3519
rect 5181 3485 5215 3519
rect 8677 3485 8711 3519
rect 8769 3485 8803 3519
rect 1869 3417 1903 3451
rect 7380 3417 7414 3451
rect 9312 3417 9346 3451
rect 3341 3349 3375 3383
rect 3801 3349 3835 3383
rect 2421 3145 2455 3179
rect 9045 3145 9079 3179
rect 9873 3145 9907 3179
rect 10241 3145 10275 3179
rect 6193 3077 6227 3111
rect 7573 3077 7607 3111
rect 2973 3009 3007 3043
rect 3525 3009 3559 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 7932 3009 7966 3043
rect 9229 3009 9263 3043
rect 10425 3009 10459 3043
rect 3157 2941 3191 2975
rect 3617 2941 3651 2975
rect 7665 2941 7699 2975
rect 7297 2873 7331 2907
rect 4721 2805 4755 2839
rect 3065 2601 3099 2635
rect 5549 2601 5583 2635
rect 8033 2601 8067 2635
rect 9781 2601 9815 2635
rect 8309 2533 8343 2567
rect 8401 2533 8435 2567
rect 3801 2465 3835 2499
rect 9505 2465 9539 2499
rect 10333 2465 10367 2499
rect 3249 2397 3283 2431
rect 7757 2397 7791 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 8953 2397 8987 2431
rect 4077 2329 4111 2363
rect 7941 2261 7975 2295
<< metal1 >>
rect 1104 11450 10764 11472
rect 1104 11398 2157 11450
rect 2209 11398 2221 11450
rect 2273 11398 2285 11450
rect 2337 11398 2349 11450
rect 2401 11398 2413 11450
rect 2465 11398 4572 11450
rect 4624 11398 4636 11450
rect 4688 11398 4700 11450
rect 4752 11398 4764 11450
rect 4816 11398 4828 11450
rect 4880 11398 6987 11450
rect 7039 11398 7051 11450
rect 7103 11398 7115 11450
rect 7167 11398 7179 11450
rect 7231 11398 7243 11450
rect 7295 11398 9402 11450
rect 9454 11398 9466 11450
rect 9518 11398 9530 11450
rect 9582 11398 9594 11450
rect 9646 11398 9658 11450
rect 9710 11398 10764 11450
rect 1104 11376 10764 11398
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 3016 11308 3249 11336
rect 3016 11296 3022 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8996 11308 9229 11336
rect 8996 11296 9002 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3142 11024 3148 11076
rect 3200 11024 3206 11076
rect 6914 11024 6920 11076
rect 6972 11024 6978 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7374 11064 7380 11076
rect 7147 11036 7380 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 9122 11024 9128 11076
rect 9180 11024 9186 11076
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3292 10968 4077 10996
rect 3292 10956 3298 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4065 10959 4123 10965
rect 7285 10999 7343 11005
rect 7285 10965 7297 10999
rect 7331 10996 7343 10999
rect 7926 10996 7932 11008
rect 7331 10968 7932 10996
rect 7331 10965 7343 10968
rect 7285 10959 7343 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 1104 10906 10923 10928
rect 1104 10854 3364 10906
rect 3416 10854 3428 10906
rect 3480 10854 3492 10906
rect 3544 10854 3556 10906
rect 3608 10854 3620 10906
rect 3672 10854 5779 10906
rect 5831 10854 5843 10906
rect 5895 10854 5907 10906
rect 5959 10854 5971 10906
rect 6023 10854 6035 10906
rect 6087 10854 8194 10906
rect 8246 10854 8258 10906
rect 8310 10854 8322 10906
rect 8374 10854 8386 10906
rect 8438 10854 8450 10906
rect 8502 10854 10609 10906
rect 10661 10854 10673 10906
rect 10725 10854 10737 10906
rect 10789 10854 10801 10906
rect 10853 10854 10865 10906
rect 10917 10854 10923 10906
rect 1104 10832 10923 10854
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 3142 10792 3148 10804
rect 2363 10764 3148 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 8110 10792 8116 10804
rect 5920 10764 8116 10792
rect 5384 10727 5442 10733
rect 5384 10693 5396 10727
rect 5430 10724 5442 10727
rect 5721 10727 5779 10733
rect 5721 10724 5733 10727
rect 5430 10696 5733 10724
rect 5430 10693 5442 10696
rect 5384 10687 5442 10693
rect 5721 10693 5733 10696
rect 5767 10693 5779 10727
rect 5721 10687 5779 10693
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 5920 10665 5948 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9122 10792 9128 10804
rect 9079 10764 9128 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 8386 10724 8392 10736
rect 6012 10696 8392 10724
rect 6012 10665 6040 10696
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 5905 10659 5963 10665
rect 3651 10628 5764 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 4430 10588 4436 10600
rect 3375 10560 4436 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5626 10548 5632 10600
rect 5684 10548 5690 10600
rect 5736 10597 5764 10628
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6972 10628 7297 10656
rect 6972 10616 6978 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7742 10656 7748 10668
rect 7607 10628 7748 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8846 10656 8852 10668
rect 8343 10628 8852 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10459 10628 10916 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7055 10560 7696 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 5736 10520 5764 10551
rect 7101 10523 7159 10529
rect 7101 10520 7113 10523
rect 5736 10492 7113 10520
rect 7101 10489 7113 10492
rect 7147 10489 7159 10523
rect 7101 10483 7159 10489
rect 7668 10464 7696 10560
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7892 10560 8033 10588
rect 7892 10548 7898 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 10888 10532 10916 10628
rect 10870 10480 10876 10532
rect 10928 10480 10934 10532
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3878 10452 3884 10464
rect 3559 10424 3884 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4246 10412 4252 10464
rect 4304 10412 4310 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 5776 10424 6377 10452
rect 5776 10412 5782 10424
rect 6365 10421 6377 10424
rect 6411 10452 6423 10455
rect 6822 10452 6828 10464
rect 6411 10424 6828 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7558 10452 7564 10464
rect 6972 10424 7564 10452
rect 6972 10412 6978 10424
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7650 10412 7656 10464
rect 7708 10412 7714 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9272 10424 10241 10452
rect 9272 10412 9278 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 1104 10362 10764 10384
rect 1104 10310 2157 10362
rect 2209 10310 2221 10362
rect 2273 10310 2285 10362
rect 2337 10310 2349 10362
rect 2401 10310 2413 10362
rect 2465 10310 4572 10362
rect 4624 10310 4636 10362
rect 4688 10310 4700 10362
rect 4752 10310 4764 10362
rect 4816 10310 4828 10362
rect 4880 10310 6987 10362
rect 7039 10310 7051 10362
rect 7103 10310 7115 10362
rect 7167 10310 7179 10362
rect 7231 10310 7243 10362
rect 7295 10310 9402 10362
rect 9454 10310 9466 10362
rect 9518 10310 9530 10362
rect 9582 10310 9594 10362
rect 9646 10310 9658 10362
rect 9710 10310 10764 10362
rect 1104 10288 10764 10310
rect 1578 10208 1584 10260
rect 1636 10208 1642 10260
rect 3234 10208 3240 10260
rect 3292 10208 3298 10260
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3476 10220 3617 10248
rect 3476 10208 3482 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 5534 10248 5540 10260
rect 3605 10211 3663 10217
rect 3804 10220 5540 10248
rect 1596 10044 1624 10208
rect 3804 10180 3832 10220
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 5718 10248 5724 10260
rect 5592 10220 5724 10248
rect 5592 10208 5598 10220
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6135 10220 7420 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 7392 10192 7420 10220
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 8202 10248 8208 10260
rect 7944 10220 8208 10248
rect 3344 10152 3832 10180
rect 3344 10121 3372 10152
rect 7374 10140 7380 10192
rect 7432 10140 7438 10192
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10081 3387 10115
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 3329 10075 3387 10081
rect 5644 10084 6285 10112
rect 5644 10056 5672 10084
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 1596 10016 2973 10044
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3694 10044 3700 10056
rect 3467 10016 3700 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 5626 10044 5632 10056
rect 3835 10016 5632 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3804 9920 3832 10007
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 3936 9948 4046 9976
rect 3936 9936 3942 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 5920 9976 5948 10007
rect 5994 10004 6000 10056
rect 6052 10004 6058 10056
rect 7668 10044 7696 10208
rect 7944 10192 7972 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8386 10208 8392 10260
rect 8444 10208 8450 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 10410 10248 10416 10260
rect 9447 10220 10416 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 7926 10140 7932 10192
rect 7984 10140 7990 10192
rect 8110 10140 8116 10192
rect 8168 10140 8174 10192
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8662 10112 8668 10124
rect 8067 10084 8668 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 6104 10016 7696 10044
rect 7929 10047 7987 10053
rect 6104 9976 6132 10016
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 7975 10016 8064 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 6546 9985 6552 9988
rect 4034 9939 4092 9945
rect 5184 9948 5764 9976
rect 5920 9948 6132 9976
rect 5184 9920 5212 9948
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 5166 9868 5172 9920
rect 5224 9868 5230 9920
rect 5258 9868 5264 9920
rect 5316 9868 5322 9920
rect 5736 9908 5764 9948
rect 6540 9939 6552 9985
rect 6546 9936 6552 9939
rect 6604 9936 6610 9988
rect 7650 9936 7656 9988
rect 7708 9936 7714 9988
rect 5994 9908 6000 9920
rect 5736 9880 6000 9908
rect 5994 9868 6000 9880
rect 6052 9908 6058 9920
rect 7668 9908 7696 9936
rect 6052 9880 7696 9908
rect 6052 9868 6058 9880
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 8036 9908 8064 10016
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 8404 10053 8432 10084
rect 8662 10072 8668 10084
rect 8720 10112 8726 10124
rect 9214 10112 9220 10124
rect 8720 10084 9220 10112
rect 8720 10072 8726 10084
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9232 10044 9260 10072
rect 9171 10016 9260 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 8588 9976 8616 10007
rect 9416 9976 9444 10211
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9631 10084 9904 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9876 10053 9904 10084
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 8588 9948 9444 9976
rect 8588 9908 8616 9948
rect 8036 9880 8616 9908
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9548 9880 9689 9908
rect 9548 9868 9554 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 1104 9818 10923 9840
rect 1104 9766 3364 9818
rect 3416 9766 3428 9818
rect 3480 9766 3492 9818
rect 3544 9766 3556 9818
rect 3608 9766 3620 9818
rect 3672 9766 5779 9818
rect 5831 9766 5843 9818
rect 5895 9766 5907 9818
rect 5959 9766 5971 9818
rect 6023 9766 6035 9818
rect 6087 9766 8194 9818
rect 8246 9766 8258 9818
rect 8310 9766 8322 9818
rect 8374 9766 8386 9818
rect 8438 9766 8450 9818
rect 8502 9766 10609 9818
rect 10661 9766 10673 9818
rect 10725 9766 10737 9818
rect 10789 9766 10801 9818
rect 10853 9766 10865 9818
rect 10917 9766 10923 9818
rect 1104 9744 10923 9766
rect 5166 9704 5172 9716
rect 4080 9676 5172 9704
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3752 9540 3893 9568
rect 3752 9528 3758 9540
rect 3881 9537 3893 9540
rect 3927 9568 3939 9571
rect 4080 9568 4108 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9664 5322 9716
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 7558 9704 7564 9716
rect 6932 9676 7564 9704
rect 3927 9540 4108 9568
rect 4157 9571 4215 9577
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 5276 9568 5304 9664
rect 6932 9636 6960 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7653 9707 7711 9713
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 8110 9704 8116 9716
rect 7699 9676 8116 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9673 8447 9707
rect 8389 9667 8447 9673
rect 5644 9608 6960 9636
rect 7208 9608 7788 9636
rect 5644 9577 5672 9608
rect 4203 9540 5304 9568
rect 5629 9571 5687 9577
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 6730 9571 6788 9577
rect 6730 9537 6742 9571
rect 6776 9568 6788 9571
rect 7208 9568 7236 9608
rect 7760 9580 7788 9608
rect 6776 9540 7236 9568
rect 6776 9537 6788 9540
rect 6730 9531 6788 9537
rect 7282 9528 7288 9580
rect 7340 9528 7346 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8404 9568 8432 9667
rect 8662 9664 8668 9716
rect 8720 9664 8726 9716
rect 8343 9540 8432 9568
rect 8573 9571 8631 9577
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 8680 9568 8708 9664
rect 9300 9639 9358 9645
rect 9300 9605 9312 9639
rect 9346 9636 9358 9639
rect 9490 9636 9496 9648
rect 9346 9608 9496 9636
rect 9346 9605 9358 9608
rect 9300 9599 9358 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 8619 9540 8708 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4488 9472 4813 9500
rect 4488 9460 4494 9472
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7484 9500 7512 9528
rect 7239 9472 7512 9500
rect 9033 9503 9091 9509
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 4246 9432 4252 9444
rect 4080 9404 4252 9432
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 4080 9373 4108 9404
rect 4246 9392 4252 9404
rect 4304 9432 4310 9444
rect 5442 9432 5448 9444
rect 4304 9404 5448 9432
rect 4304 9392 4310 9404
rect 5442 9392 5448 9404
rect 5500 9432 5506 9444
rect 6840 9432 6868 9460
rect 9048 9432 9076 9463
rect 5500 9404 6316 9432
rect 6840 9404 9076 9432
rect 5500 9392 5506 9404
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6052 9336 6193 9364
rect 6052 9324 6058 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6288 9364 6316 9404
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6288 9336 7297 9364
rect 6181 9327 6239 9333
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7926 9364 7932 9376
rect 7432 9336 7932 9364
rect 7432 9324 7438 9336
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8110 9324 8116 9376
rect 8168 9324 8174 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10459 9336 10824 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 1104 9274 10764 9296
rect 1104 9222 2157 9274
rect 2209 9222 2221 9274
rect 2273 9222 2285 9274
rect 2337 9222 2349 9274
rect 2401 9222 2413 9274
rect 2465 9222 4572 9274
rect 4624 9222 4636 9274
rect 4688 9222 4700 9274
rect 4752 9222 4764 9274
rect 4816 9222 4828 9274
rect 4880 9222 6987 9274
rect 7039 9222 7051 9274
rect 7103 9222 7115 9274
rect 7167 9222 7179 9274
rect 7231 9222 7243 9274
rect 7295 9222 9402 9274
rect 9454 9222 9466 9274
rect 9518 9222 9530 9274
rect 9582 9222 9594 9274
rect 9646 9222 9658 9274
rect 9710 9222 10764 9274
rect 1104 9200 10764 9222
rect 3602 9120 3608 9172
rect 3660 9120 3666 9172
rect 4430 9120 4436 9172
rect 4488 9120 4494 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5074 9160 5080 9172
rect 4939 9132 5080 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5534 9120 5540 9172
rect 5592 9120 5598 9172
rect 3620 9024 3648 9120
rect 4448 9092 4476 9120
rect 6730 9092 6736 9104
rect 4448 9064 6736 9092
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 3620 8996 4261 9024
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 5442 8984 5448 9036
rect 5500 8984 5506 9036
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 5460 8956 5488 8984
rect 5399 8928 5488 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6196 8965 6224 9064
rect 6730 9052 6736 9064
rect 6788 9092 6794 9104
rect 7834 9092 7840 9104
rect 6788 9064 7840 9092
rect 6788 9052 6794 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10796 9024 10824 9336
rect 10459 8996 10824 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9723 8928 9781 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6365 8891 6423 8897
rect 6365 8888 6377 8891
rect 5684 8860 6377 8888
rect 5684 8848 5690 8860
rect 6365 8857 6377 8860
rect 6411 8857 6423 8891
rect 6365 8851 6423 8857
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7558 8888 7564 8900
rect 7340 8860 7564 8888
rect 7340 8848 7346 8860
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 7653 8891 7711 8897
rect 7653 8857 7665 8891
rect 7699 8888 7711 8891
rect 7742 8888 7748 8900
rect 7699 8860 7748 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 7742 8848 7748 8860
rect 7800 8848 7806 8900
rect 7837 8891 7895 8897
rect 7837 8857 7849 8891
rect 7883 8888 7895 8891
rect 7926 8888 7932 8900
rect 7883 8860 7932 8888
rect 7883 8857 7895 8860
rect 7837 8851 7895 8857
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 9858 8888 9864 8900
rect 8076 8860 9864 8888
rect 8076 8848 8082 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 7300 8820 7328 8848
rect 5859 8792 7328 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 9214 8780 9220 8832
rect 9272 8820 9278 8832
rect 9585 8823 9643 8829
rect 9585 8820 9597 8823
rect 9272 8792 9597 8820
rect 9272 8780 9278 8792
rect 9585 8789 9597 8792
rect 9631 8789 9643 8823
rect 9585 8783 9643 8789
rect 1104 8730 10923 8752
rect 1104 8678 3364 8730
rect 3416 8678 3428 8730
rect 3480 8678 3492 8730
rect 3544 8678 3556 8730
rect 3608 8678 3620 8730
rect 3672 8678 5779 8730
rect 5831 8678 5843 8730
rect 5895 8678 5907 8730
rect 5959 8678 5971 8730
rect 6023 8678 6035 8730
rect 6087 8678 8194 8730
rect 8246 8678 8258 8730
rect 8310 8678 8322 8730
rect 8374 8678 8386 8730
rect 8438 8678 8450 8730
rect 8502 8678 10609 8730
rect 10661 8678 10673 8730
rect 10725 8678 10737 8730
rect 10789 8678 10801 8730
rect 10853 8678 10865 8730
rect 10917 8678 10923 8730
rect 1104 8656 10923 8678
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 6564 8588 7481 8616
rect 6564 8557 6592 8588
rect 7469 8585 7481 8588
rect 7515 8616 7527 8619
rect 7650 8616 7656 8628
rect 7515 8588 7656 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 8018 8576 8024 8628
rect 8076 8576 8082 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 6549 8551 6607 8557
rect 6549 8517 6561 8551
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 6779 8520 7328 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 7300 8492 7328 8520
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 3694 8480 3700 8492
rect 2990 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3988 8452 4077 8480
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 3988 8356 4016 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 8036 8480 8064 8576
rect 7607 8452 8064 8480
rect 8128 8480 8156 8576
rect 8185 8483 8243 8489
rect 8185 8480 8197 8483
rect 8128 8452 8197 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 8185 8449 8197 8452
rect 8231 8449 8243 8483
rect 8185 8443 8243 8449
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6822 8412 6828 8424
rect 6420 8384 6828 8412
rect 6420 8372 6426 8384
rect 6822 8372 6828 8384
rect 6880 8412 6886 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 6880 8384 7941 8412
rect 6880 8372 6886 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 3970 8344 3976 8356
rect 3375 8316 3976 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7834 8344 7840 8356
rect 7147 8316 7840 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 3878 8236 3884 8288
rect 3936 8236 3942 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 5592 8248 6377 8276
rect 5592 8236 5598 8248
rect 6365 8245 6377 8248
rect 6411 8276 6423 8279
rect 6822 8276 6828 8288
rect 6411 8248 6828 8276
rect 6411 8245 6423 8248
rect 6365 8239 6423 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 1104 8186 10764 8208
rect 1104 8134 2157 8186
rect 2209 8134 2221 8186
rect 2273 8134 2285 8186
rect 2337 8134 2349 8186
rect 2401 8134 2413 8186
rect 2465 8134 4572 8186
rect 4624 8134 4636 8186
rect 4688 8134 4700 8186
rect 4752 8134 4764 8186
rect 4816 8134 4828 8186
rect 4880 8134 6987 8186
rect 7039 8134 7051 8186
rect 7103 8134 7115 8186
rect 7167 8134 7179 8186
rect 7231 8134 7243 8186
rect 7295 8134 9402 8186
rect 9454 8134 9466 8186
rect 9518 8134 9530 8186
rect 9582 8134 9594 8186
rect 9646 8134 9658 8186
rect 9710 8134 10764 8186
rect 1104 8112 10764 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1854 8072 1860 8084
rect 1627 8044 1860 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7466 8072 7472 8084
rect 7147 8044 7472 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 9858 8032 9864 8084
rect 9916 8032 9922 8084
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 9122 8004 9128 8016
rect 6880 7976 9128 8004
rect 6880 7964 6886 7976
rect 9122 7964 9128 7976
rect 9180 8004 9186 8016
rect 9180 7976 9536 8004
rect 9180 7964 9186 7976
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 2866 7936 2872 7948
rect 2087 7908 2872 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 3016 7908 3065 7936
rect 3016 7896 3022 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3053 7899 3111 7905
rect 3344 7908 3525 7936
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 3344 7868 3372 7908
rect 3513 7905 3525 7908
rect 3559 7936 3571 7939
rect 3878 7936 3884 7948
rect 3559 7908 3884 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 9508 7945 9536 7976
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 1995 7840 3372 7868
rect 3421 7871 3479 7877
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 3436 7800 3464 7831
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 3292 7772 3464 7800
rect 5261 7803 5319 7809
rect 3292 7760 3298 7772
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 6178 7800 6184 7812
rect 5307 7772 6184 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 9784 7800 9812 7831
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10275 7840 10364 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10060 7800 10088 7831
rect 9784 7772 9996 7800
rect 10060 7772 10272 7800
rect 9968 7744 9996 7772
rect 10244 7744 10272 7772
rect 10336 7744 10364 7840
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 6362 7732 6368 7744
rect 3844 7704 6368 7732
rect 3844 7692 3850 7704
rect 6362 7692 6368 7704
rect 6420 7732 6426 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6420 7704 6561 7732
rect 6420 7692 6426 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 7926 7692 7932 7744
rect 7984 7692 7990 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9766 7732 9772 7744
rect 9447 7704 9772 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 9950 7692 9956 7744
rect 10008 7692 10014 7744
rect 10134 7692 10140 7744
rect 10192 7692 10198 7744
rect 10226 7692 10232 7744
rect 10284 7692 10290 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 1104 7642 10923 7664
rect 1104 7590 3364 7642
rect 3416 7590 3428 7642
rect 3480 7590 3492 7642
rect 3544 7590 3556 7642
rect 3608 7590 3620 7642
rect 3672 7590 5779 7642
rect 5831 7590 5843 7642
rect 5895 7590 5907 7642
rect 5959 7590 5971 7642
rect 6023 7590 6035 7642
rect 6087 7590 8194 7642
rect 8246 7590 8258 7642
rect 8310 7590 8322 7642
rect 8374 7590 8386 7642
rect 8438 7590 8450 7642
rect 8502 7590 10609 7642
rect 10661 7590 10673 7642
rect 10725 7590 10737 7642
rect 10789 7590 10801 7642
rect 10853 7590 10865 7642
rect 10917 7590 10923 7642
rect 1104 7568 10923 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 3786 7528 3792 7540
rect 1636 7500 3792 7528
rect 1636 7488 1642 7500
rect 1688 7401 1716 7500
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 3602 7392 3608 7404
rect 3082 7364 3608 7392
rect 1673 7355 1731 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3712 7392 3740 7500
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 7466 7528 7472 7540
rect 6472 7500 7472 7528
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6472 7460 6500 7500
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 8665 7531 8723 7537
rect 8665 7528 8677 7531
rect 8628 7500 8677 7528
rect 8628 7488 8634 7500
rect 8665 7497 8677 7500
rect 8711 7497 8723 7531
rect 8665 7491 8723 7497
rect 8938 7488 8944 7540
rect 8996 7488 9002 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 9272 7500 9505 7528
rect 9272 7488 9278 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 9493 7491 9551 7497
rect 5592 7432 5948 7460
rect 5592 7420 5598 7432
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3712 7364 3801 7392
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 5626 7392 5632 7404
rect 5198 7378 5632 7392
rect 3789 7355 3847 7361
rect 5184 7364 5632 7378
rect 1946 7284 1952 7336
rect 2004 7284 2010 7336
rect 2958 7284 2964 7336
rect 3016 7284 3022 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3804 7296 4077 7324
rect 2976 7256 3004 7284
rect 3804 7256 3832 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 2976 7228 3832 7256
rect 3418 7148 3424 7200
rect 3476 7148 3482 7200
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 5184 7188 5212 7364
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5920 7401 5948 7432
rect 6196 7432 6500 7460
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 6196 7333 6224 7432
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8297 7463 8355 7469
rect 8297 7429 8309 7463
rect 8343 7460 8355 7463
rect 8956 7460 8984 7488
rect 8343 7432 8984 7460
rect 8343 7429 8355 7432
rect 8297 7423 8355 7429
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 6472 7364 6633 7392
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7293 6239 7327
rect 6472 7324 6500 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 8036 7392 8064 7420
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8036 7364 8769 7392
rect 6621 7355 6679 7361
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 6181 7287 6239 7293
rect 6380 7296 6500 7324
rect 5721 7259 5779 7265
rect 5721 7225 5733 7259
rect 5767 7256 5779 7259
rect 6380 7256 6408 7296
rect 7834 7284 7840 7336
rect 7892 7324 7898 7336
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7892 7296 8033 7324
rect 7892 7284 7898 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 8570 7324 8576 7336
rect 8251 7296 8576 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 5767 7228 6408 7256
rect 8036 7256 8064 7287
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8662 7256 8668 7268
rect 8036 7228 8668 7256
rect 5767 7225 5779 7228
rect 5721 7219 5779 7225
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 8956 7256 8984 7355
rect 9140 7324 9168 7488
rect 10318 7460 10324 7472
rect 9324 7432 10324 7460
rect 9324 7404 9352 7432
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9447 7364 10149 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 10137 7361 10149 7364
rect 10183 7392 10195 7395
rect 10226 7392 10232 7404
rect 10183 7364 10232 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9140 7296 9229 7324
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 8956 7228 9996 7256
rect 9968 7200 9996 7228
rect 3660 7160 5212 7188
rect 3660 7148 3666 7160
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 6135 7160 8953 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 8941 7157 8953 7160
rect 8987 7157 8999 7191
rect 8941 7151 8999 7157
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 1104 7098 10764 7120
rect 1104 7046 2157 7098
rect 2209 7046 2221 7098
rect 2273 7046 2285 7098
rect 2337 7046 2349 7098
rect 2401 7046 2413 7098
rect 2465 7046 4572 7098
rect 4624 7046 4636 7098
rect 4688 7046 4700 7098
rect 4752 7046 4764 7098
rect 4816 7046 4828 7098
rect 4880 7046 6987 7098
rect 7039 7046 7051 7098
rect 7103 7046 7115 7098
rect 7167 7046 7179 7098
rect 7231 7046 7243 7098
rect 7295 7046 9402 7098
rect 9454 7046 9466 7098
rect 9518 7046 9530 7098
rect 9582 7046 9594 7098
rect 9646 7046 9658 7098
rect 9710 7046 10764 7098
rect 1104 7024 10764 7046
rect 1946 6944 1952 6996
rect 2004 6944 2010 6996
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3878 6984 3884 6996
rect 2924 6956 3884 6984
rect 2924 6944 2930 6956
rect 3878 6944 3884 6956
rect 3936 6984 3942 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 3936 6956 3985 6984
rect 3936 6944 3942 6956
rect 3973 6953 3985 6956
rect 4019 6953 4031 6987
rect 3973 6947 4031 6953
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 9306 6916 9312 6928
rect 8803 6888 9312 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 9306 6876 9312 6888
rect 9364 6916 9370 6928
rect 9364 6888 9536 6916
rect 9364 6876 9370 6888
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 1912 6820 2145 6848
rect 1912 6808 1918 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 2133 6811 2191 6817
rect 3252 6820 4997 6848
rect 3252 6792 3280 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5534 6848 5540 6860
rect 5307 6820 5540 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 9508 6857 9536 6888
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 9916 6820 10241 6848
rect 9916 6808 9922 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2958 6780 2964 6792
rect 2271 6752 2964 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7423 6752 8616 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 3418 6712 3424 6724
rect 2792 6684 3424 6712
rect 2792 6656 2820 6684
rect 3418 6672 3424 6684
rect 3476 6712 3482 6724
rect 3804 6712 3832 6743
rect 3476 6684 3832 6712
rect 3476 6672 3482 6684
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4212 6684 5365 6712
rect 4212 6672 4218 6684
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 7644 6715 7702 6721
rect 7644 6681 7656 6715
rect 7690 6712 7702 6715
rect 7742 6712 7748 6724
rect 7690 6684 7748 6712
rect 7690 6681 7702 6684
rect 7644 6675 7702 6681
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 8588 6656 8616 6752
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6236 6616 6653 6644
rect 6236 6604 6242 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 8904 6616 9689 6644
rect 8904 6604 8910 6616
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 1104 6554 10923 6576
rect 1104 6502 3364 6554
rect 3416 6502 3428 6554
rect 3480 6502 3492 6554
rect 3544 6502 3556 6554
rect 3608 6502 3620 6554
rect 3672 6502 5779 6554
rect 5831 6502 5843 6554
rect 5895 6502 5907 6554
rect 5959 6502 5971 6554
rect 6023 6502 6035 6554
rect 6087 6502 8194 6554
rect 8246 6502 8258 6554
rect 8310 6502 8322 6554
rect 8374 6502 8386 6554
rect 8438 6502 8450 6554
rect 8502 6502 10609 6554
rect 10661 6502 10673 6554
rect 10725 6502 10737 6554
rect 10789 6502 10801 6554
rect 10853 6502 10865 6554
rect 10917 6502 10923 6554
rect 1104 6480 10923 6502
rect 7742 6400 7748 6452
rect 7800 6400 7806 6452
rect 7926 6400 7932 6452
rect 7984 6400 7990 6452
rect 8846 6400 8852 6452
rect 8904 6400 8910 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 5258 6304 5264 6316
rect 4663 6276 5264 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 7944 6313 7972 6400
rect 8864 6372 8892 6400
rect 8496 6344 8892 6372
rect 8956 6372 8984 6403
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10284 6412 10425 6440
rect 10284 6400 10290 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 9278 6375 9336 6381
rect 9278 6372 9290 6375
rect 8956 6344 9290 6372
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5684 6276 6377 6304
rect 5684 6264 5690 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 3234 6196 3240 6248
rect 3292 6196 3298 6248
rect 3878 6196 3884 6248
rect 3936 6196 3942 6248
rect 8496 6245 8524 6344
rect 9278 6341 9290 6344
rect 9324 6341 9336 6375
rect 9278 6335 9336 6341
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8662 6304 8668 6316
rect 8619 6276 8668 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4172 6208 4537 6236
rect 3252 6168 3280 6196
rect 4172 6168 4200 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8481 6199 8539 6205
rect 8588 6208 9045 6236
rect 3252 6140 4200 6168
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 5092 6168 5120 6199
rect 4387 6140 5120 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 8588 6112 8616 6208
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5534 6100 5540 6112
rect 5031 6072 5540 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 6328 6072 6561 6100
rect 6328 6060 6334 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 1104 6010 10764 6032
rect 1104 5958 2157 6010
rect 2209 5958 2221 6010
rect 2273 5958 2285 6010
rect 2337 5958 2349 6010
rect 2401 5958 2413 6010
rect 2465 5958 4572 6010
rect 4624 5958 4636 6010
rect 4688 5958 4700 6010
rect 4752 5958 4764 6010
rect 4816 5958 4828 6010
rect 4880 5958 6987 6010
rect 7039 5958 7051 6010
rect 7103 5958 7115 6010
rect 7167 5958 7179 6010
rect 7231 5958 7243 6010
rect 7295 5958 9402 6010
rect 9454 5958 9466 6010
rect 9518 5958 9530 6010
rect 9582 5958 9594 6010
rect 9646 5958 9658 6010
rect 9710 5958 10764 6010
rect 1104 5936 10764 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 7650 5896 7656 5908
rect 7331 5868 7656 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 7650 5856 7656 5868
rect 7708 5896 7714 5908
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 7708 5868 8401 5896
rect 7708 5856 7714 5868
rect 8389 5865 8401 5868
rect 8435 5896 8447 5899
rect 8846 5896 8852 5908
rect 8435 5868 8852 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9824 5868 10057 5896
rect 9824 5856 9830 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5797 2467 5831
rect 2409 5791 2467 5797
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2424 5760 2452 5791
rect 2271 5732 2452 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2866 5720 2872 5772
rect 2924 5720 2930 5772
rect 3252 5760 3280 5856
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 3252 5732 3341 5760
rect 3329 5729 3341 5732
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3605 5763 3663 5769
rect 3605 5729 3617 5763
rect 3651 5760 3663 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3651 5732 4077 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2179 5664 2268 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2240 5568 2268 5664
rect 2774 5652 2780 5704
rect 2832 5652 2838 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3970 5692 3976 5704
rect 3283 5664 3976 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3970 5652 3976 5664
rect 4028 5692 4034 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4028 5664 5457 5692
rect 4028 5652 4034 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 8711 5664 9076 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 5552 5624 5580 5655
rect 5552 5596 5672 5624
rect 5644 5568 5672 5596
rect 6270 5584 6276 5636
rect 6328 5584 6334 5636
rect 9048 5568 9076 5664
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 2222 5516 2228 5568
rect 2280 5516 2286 5568
rect 4706 5516 4712 5568
rect 4764 5516 4770 5568
rect 5258 5516 5264 5568
rect 5316 5516 5322 5568
rect 5626 5516 5632 5568
rect 5684 5516 5690 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7892 5528 8217 5556
rect 7892 5516 7898 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 9030 5516 9036 5568
rect 9088 5516 9094 5568
rect 9214 5516 9220 5568
rect 9272 5516 9278 5568
rect 1104 5466 10923 5488
rect 1104 5414 3364 5466
rect 3416 5414 3428 5466
rect 3480 5414 3492 5466
rect 3544 5414 3556 5466
rect 3608 5414 3620 5466
rect 3672 5414 5779 5466
rect 5831 5414 5843 5466
rect 5895 5414 5907 5466
rect 5959 5414 5971 5466
rect 6023 5414 6035 5466
rect 6087 5414 8194 5466
rect 8246 5414 8258 5466
rect 8310 5414 8322 5466
rect 8374 5414 8386 5466
rect 8438 5414 8450 5466
rect 8502 5414 10609 5466
rect 10661 5414 10673 5466
rect 10725 5414 10737 5466
rect 10789 5414 10801 5466
rect 10853 5414 10865 5466
rect 10917 5414 10923 5466
rect 1104 5392 10923 5414
rect 3970 5312 3976 5364
rect 4028 5312 4034 5364
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 4764 5324 5488 5352
rect 4764 5312 4770 5324
rect 5460 5293 5488 5324
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6328 5324 6776 5352
rect 6328 5312 6334 5324
rect 5445 5287 5503 5293
rect 5445 5253 5457 5287
rect 5491 5253 5503 5287
rect 5445 5247 5503 5253
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 5592 5256 6653 5284
rect 5592 5244 5598 5256
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 6748 5284 6776 5324
rect 8748 5287 8806 5293
rect 6748 5256 7130 5284
rect 6641 5247 6699 5253
rect 8748 5253 8760 5287
rect 8794 5284 8806 5287
rect 9214 5284 9220 5296
rect 8794 5256 9220 5284
rect 8794 5253 8806 5256
rect 8748 5247 8806 5253
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 8481 5219 8539 5225
rect 1946 5108 1952 5160
rect 2004 5108 2010 5160
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 2682 5148 2688 5160
rect 2280 5120 2688 5148
rect 2280 5108 2286 5120
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3344 5148 3372 5202
rect 4356 5148 4384 5202
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 8570 5216 8576 5228
rect 8527 5188 8576 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 3292 5120 4384 5148
rect 5644 5120 5733 5148
rect 3292 5108 3298 5120
rect 5644 5024 5672 5120
rect 5721 5117 5733 5120
rect 5767 5148 5779 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5767 5120 6377 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 3694 4972 3700 5024
rect 3752 4972 3758 5024
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8754 5012 8760 5024
rect 8159 4984 8760 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8754 4972 8760 4984
rect 8812 5012 8818 5024
rect 9122 5012 9128 5024
rect 8812 4984 9128 5012
rect 8812 4972 8818 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9858 4972 9864 5024
rect 9916 4972 9922 5024
rect 1104 4922 10764 4944
rect 1104 4870 2157 4922
rect 2209 4870 2221 4922
rect 2273 4870 2285 4922
rect 2337 4870 2349 4922
rect 2401 4870 2413 4922
rect 2465 4870 4572 4922
rect 4624 4870 4636 4922
rect 4688 4870 4700 4922
rect 4752 4870 4764 4922
rect 4816 4870 4828 4922
rect 4880 4870 6987 4922
rect 7039 4870 7051 4922
rect 7103 4870 7115 4922
rect 7167 4870 7179 4922
rect 7231 4870 7243 4922
rect 7295 4870 9402 4922
rect 9454 4870 9466 4922
rect 9518 4870 9530 4922
rect 9582 4870 9594 4922
rect 9646 4870 9658 4922
rect 9710 4870 10764 4922
rect 1104 4848 10764 4870
rect 3694 4768 3700 4820
rect 3752 4768 3758 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8312 4780 9321 4808
rect 3712 4672 3740 4768
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 8312 4740 8340 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9766 4808 9772 4820
rect 9723 4780 9772 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 7616 4712 8340 4740
rect 7616 4700 7622 4712
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 9217 4743 9275 4749
rect 9217 4740 9229 4743
rect 8904 4712 9229 4740
rect 8904 4700 8910 4712
rect 9217 4709 9229 4712
rect 9263 4709 9275 4743
rect 9217 4703 9275 4709
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 3712 4644 4169 4672
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 8662 4632 8668 4684
rect 8720 4632 8726 4684
rect 9122 4632 9128 4684
rect 9180 4632 9186 4684
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9916 4644 10333 4672
rect 9916 4632 9922 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4448 4480 4476 4567
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9030 4604 9036 4616
rect 8987 4576 9036 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9030 4564 9036 4576
rect 9088 4604 9094 4616
rect 9214 4604 9220 4616
rect 9088 4576 9220 4604
rect 9088 4564 9094 4576
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9447 4576 9781 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 7926 4428 7932 4480
rect 7984 4428 7990 4480
rect 8018 4428 8024 4480
rect 8076 4428 8082 4480
rect 1104 4378 10923 4400
rect 1104 4326 3364 4378
rect 3416 4326 3428 4378
rect 3480 4326 3492 4378
rect 3544 4326 3556 4378
rect 3608 4326 3620 4378
rect 3672 4326 5779 4378
rect 5831 4326 5843 4378
rect 5895 4326 5907 4378
rect 5959 4326 5971 4378
rect 6023 4326 6035 4378
rect 6087 4326 8194 4378
rect 8246 4326 8258 4378
rect 8310 4326 8322 4378
rect 8374 4326 8386 4378
rect 8438 4326 8450 4378
rect 8502 4326 10609 4378
rect 10661 4326 10673 4378
rect 10725 4326 10737 4378
rect 10789 4326 10801 4378
rect 10853 4326 10865 4378
rect 10917 4326 10923 4378
rect 1104 4304 10923 4326
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 7282 4264 7288 4276
rect 7239 4236 7288 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8159 4236 9996 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 7944 4168 8156 4196
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 3436 4100 4169 4128
rect 3436 4069 3464 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 5534 4128 5540 4140
rect 4663 4100 5540 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 3970 4060 3976 4072
rect 3743 4032 3976 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4172 4060 4200 4091
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 4430 4060 4436 4072
rect 4172 4032 4436 4060
rect 4065 4023 4123 4029
rect 4080 3992 4108 4023
rect 4430 4020 4436 4032
rect 4488 4060 4494 4072
rect 4525 4063 4583 4069
rect 4525 4060 4537 4063
rect 4488 4032 4537 4060
rect 4488 4020 4494 4032
rect 4525 4029 4537 4032
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4060 5043 4063
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5031 4032 5181 4060
rect 5031 4029 5043 4032
rect 4985 4023 5043 4029
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 7484 4060 7512 4091
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 7944 4137 7972 4168
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7800 4100 7941 4128
rect 7800 4088 7806 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 8036 4060 8064 4088
rect 7484 4032 8064 4060
rect 8128 4060 8156 4168
rect 8754 4088 8760 4140
rect 8812 4088 8818 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 9858 4128 9864 4140
rect 9815 4100 9864 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9968 4128 9996 4236
rect 10042 4128 10048 4140
rect 9968 4100 10048 4128
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 8128 4032 8340 4060
rect 5169 4023 5227 4029
rect 5258 3992 5264 4004
rect 2746 3964 3832 3992
rect 4080 3964 5264 3992
rect 2746 3936 2774 3964
rect 2682 3884 2688 3936
rect 2740 3896 2774 3936
rect 3804 3933 3832 3964
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 8202 3992 8208 4004
rect 7791 3964 8208 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 3789 3927 3847 3933
rect 2740 3884 2746 3896
rect 3789 3893 3801 3927
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5776 3896 5825 3924
rect 5776 3884 5782 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 8312 3924 8340 4032
rect 8846 4020 8852 4072
rect 8904 4069 8910 4072
rect 8904 4063 8953 4069
rect 8904 4029 8907 4063
rect 8941 4029 8953 4063
rect 8904 4023 8953 4029
rect 8904 4020 8910 4023
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9950 4020 9956 4072
rect 10008 4020 10014 4072
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9214 3924 9220 3936
rect 8312 3896 9220 3924
rect 5813 3887 5871 3893
rect 9214 3884 9220 3896
rect 9272 3924 9278 3936
rect 9324 3924 9352 3955
rect 9272 3896 9352 3924
rect 9272 3884 9278 3896
rect 1104 3834 10764 3856
rect 1104 3782 2157 3834
rect 2209 3782 2221 3834
rect 2273 3782 2285 3834
rect 2337 3782 2349 3834
rect 2401 3782 2413 3834
rect 2465 3782 4572 3834
rect 4624 3782 4636 3834
rect 4688 3782 4700 3834
rect 4752 3782 4764 3834
rect 4816 3782 4828 3834
rect 4880 3782 6987 3834
rect 7039 3782 7051 3834
rect 7103 3782 7115 3834
rect 7167 3782 7179 3834
rect 7231 3782 7243 3834
rect 7295 3782 9402 3834
rect 9454 3782 9466 3834
rect 9518 3782 9530 3834
rect 9582 3782 9594 3834
rect 9646 3782 9658 3834
rect 9710 3782 10764 3834
rect 1104 3760 10764 3782
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3384 3692 4537 3720
rect 3384 3680 3390 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 5524 3723 5582 3729
rect 5524 3689 5536 3723
rect 5570 3720 5582 3723
rect 5718 3720 5724 3732
rect 5570 3692 5724 3720
rect 5570 3689 5582 3692
rect 5524 3683 5582 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7742 3720 7748 3732
rect 7055 3692 7748 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8662 3720 8668 3732
rect 8527 3692 8668 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10318 3720 10324 3732
rect 10008 3692 10324 3720
rect 10008 3680 10014 3692
rect 10318 3680 10324 3692
rect 10376 3720 10382 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 10376 3692 10425 3720
rect 10376 3680 10382 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1946 3584 1952 3596
rect 1627 3556 1952 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1946 3544 1952 3556
rect 2004 3584 2010 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 2004 3556 5273 3584
rect 2004 3544 2010 3556
rect 3712 3528 3740 3556
rect 5261 3553 5273 3556
rect 5307 3584 5319 3587
rect 5626 3584 5632 3596
rect 5307 3556 5632 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5626 3544 5632 3556
rect 5684 3584 5690 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 5684 3556 7113 3584
rect 5684 3544 5690 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 8570 3584 8576 3596
rect 7101 3547 7159 3553
rect 8128 3556 8576 3584
rect 3234 3516 3240 3528
rect 2990 3488 3240 3516
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3694 3476 3700 3528
rect 3752 3476 3758 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 7116 3516 7144 3547
rect 8128 3516 8156 3556
rect 8570 3544 8576 3556
rect 8628 3584 8634 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8628 3556 9045 3584
rect 8628 3544 8634 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 7116 3488 8156 3516
rect 1854 3408 1860 3460
rect 1912 3408 1918 3460
rect 4356 3448 4384 3479
rect 3344 3420 4384 3448
rect 3344 3389 3372 3420
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3349 3387 3383
rect 3329 3343 3387 3349
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 5184 3380 5212 3479
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 5500 3420 6026 3448
rect 5500 3408 5506 3420
rect 5534 3380 5540 3392
rect 5184 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5920 3380 5948 3420
rect 6270 3380 6276 3392
rect 5920 3352 6276 3380
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7116 3380 7144 3488
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8260 3488 8677 3516
rect 8260 3476 8266 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 9122 3516 9128 3528
rect 8803 3488 9128 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 7368 3451 7426 3457
rect 7368 3417 7380 3451
rect 7414 3448 7426 3451
rect 7926 3448 7932 3460
rect 7414 3420 7932 3448
rect 7414 3417 7426 3420
rect 7368 3411 7426 3417
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 7282 3380 7288 3392
rect 7116 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 8772 3380 8800 3479
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9300 3451 9358 3457
rect 9300 3417 9312 3451
rect 9346 3448 9358 3451
rect 9858 3448 9864 3460
rect 9346 3420 9864 3448
rect 9346 3417 9358 3420
rect 9300 3411 9358 3417
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 7800 3352 8800 3380
rect 7800 3340 7806 3352
rect 1104 3290 10923 3312
rect 1104 3238 3364 3290
rect 3416 3238 3428 3290
rect 3480 3238 3492 3290
rect 3544 3238 3556 3290
rect 3608 3238 3620 3290
rect 3672 3238 5779 3290
rect 5831 3238 5843 3290
rect 5895 3238 5907 3290
rect 5959 3238 5971 3290
rect 6023 3238 6035 3290
rect 6087 3238 8194 3290
rect 8246 3238 8258 3290
rect 8310 3238 8322 3290
rect 8374 3238 8386 3290
rect 8438 3238 8450 3290
rect 8502 3238 10609 3290
rect 10661 3238 10673 3290
rect 10725 3238 10737 3290
rect 10789 3238 10801 3290
rect 10853 3238 10865 3290
rect 10917 3238 10923 3290
rect 1104 3216 10923 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 2409 3179 2467 3185
rect 2409 3176 2421 3179
rect 1912 3148 2421 3176
rect 1912 3136 1918 3148
rect 2409 3145 2421 3148
rect 2455 3145 2467 3179
rect 2409 3139 2467 3145
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 7834 3176 7840 3188
rect 7208 3148 7840 3176
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2924 3012 2973 3040
rect 2924 3000 2930 3012
rect 2961 3009 2973 3012
rect 3007 3040 3019 3043
rect 3513 3043 3571 3049
rect 3007 3012 3188 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3160 2981 3188 3012
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3804 3040 3832 3136
rect 6178 3068 6184 3120
rect 6236 3068 6242 3120
rect 7208 3049 7236 3148
rect 7834 3136 7840 3148
rect 7892 3176 7898 3188
rect 8386 3176 8392 3188
rect 7892 3148 8392 3176
rect 7892 3136 7898 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9030 3136 9036 3188
rect 9088 3136 9094 3188
rect 9858 3136 9864 3188
rect 9916 3136 9922 3188
rect 10229 3179 10287 3185
rect 10229 3145 10241 3179
rect 10275 3176 10287 3179
rect 10410 3176 10416 3188
rect 10275 3148 10416 3176
rect 10275 3145 10287 3148
rect 10229 3139 10287 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 7561 3111 7619 3117
rect 7561 3077 7573 3111
rect 7607 3108 7619 3111
rect 7607 3080 9260 3108
rect 7607 3077 7619 3080
rect 7561 3071 7619 3077
rect 3559 3012 3832 3040
rect 7101 3043 7159 3049
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 5534 2972 5540 2984
rect 3651 2944 5540 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 4062 2904 4068 2916
rect 3292 2876 4068 2904
rect 3292 2864 3298 2876
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 3752 2808 4721 2836
rect 3752 2796 3758 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 7116 2836 7144 3003
rect 7300 2972 7328 3068
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7742 3040 7748 3052
rect 7423 3012 7748 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7926 3049 7932 3052
rect 7920 3003 7932 3049
rect 7926 3000 7932 3003
rect 7984 3000 7990 3052
rect 9232 3049 9260 3080
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3040 10471 3043
rect 10870 3040 10876 3052
rect 10459 3012 10876 3040
rect 10459 3009 10471 3012
rect 10413 3003 10471 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7300 2944 7665 2972
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 7558 2904 7564 2916
rect 7331 2876 7564 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 9766 2836 9772 2848
rect 7116 2808 9772 2836
rect 4709 2799 4767 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 1104 2746 10764 2768
rect 1104 2694 2157 2746
rect 2209 2694 2221 2746
rect 2273 2694 2285 2746
rect 2337 2694 2349 2746
rect 2401 2694 2413 2746
rect 2465 2694 4572 2746
rect 4624 2694 4636 2746
rect 4688 2694 4700 2746
rect 4752 2694 4764 2746
rect 4816 2694 4828 2746
rect 4880 2694 6987 2746
rect 7039 2694 7051 2746
rect 7103 2694 7115 2746
rect 7167 2694 7179 2746
rect 7231 2694 7243 2746
rect 7295 2694 9402 2746
rect 9454 2694 9466 2746
rect 9518 2694 9530 2746
rect 9582 2694 9594 2746
rect 9646 2694 9658 2746
rect 9710 2694 10764 2746
rect 1104 2672 10764 2694
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 2924 2604 3065 2632
rect 2924 2592 2930 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 7558 2592 7564 2644
rect 7616 2592 7622 2644
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7984 2604 8033 2632
rect 7984 2592 7990 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8021 2595 8079 2601
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 7576 2564 7604 2592
rect 8297 2567 8355 2573
rect 8297 2564 8309 2567
rect 7576 2536 8309 2564
rect 8297 2533 8309 2536
rect 8343 2533 8355 2567
rect 8297 2527 8355 2533
rect 8386 2524 8392 2576
rect 8444 2524 8450 2576
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3752 2468 3801 2496
rect 3752 2456 3758 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9088 2468 9505 2496
rect 9088 2456 9094 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 10318 2456 10324 2508
rect 10376 2456 10382 2508
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3016 2400 3249 2428
rect 3016 2388 3022 2400
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 4028 2332 4077 2360
rect 4028 2320 4034 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 4065 2323 4123 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 7760 2360 7788 2391
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 8168 2400 8217 2428
rect 8168 2388 8174 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8527 2400 8953 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 8754 2360 8760 2372
rect 4212 2332 4554 2360
rect 7760 2332 8760 2360
rect 4212 2320 4218 2332
rect 4448 2292 4476 2332
rect 8754 2320 8760 2332
rect 8812 2320 8818 2372
rect 5442 2292 5448 2304
rect 4448 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 7929 2295 7987 2301
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8938 2292 8944 2304
rect 7975 2264 8944 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 1104 2202 10923 2224
rect 1104 2150 3364 2202
rect 3416 2150 3428 2202
rect 3480 2150 3492 2202
rect 3544 2150 3556 2202
rect 3608 2150 3620 2202
rect 3672 2150 5779 2202
rect 5831 2150 5843 2202
rect 5895 2150 5907 2202
rect 5959 2150 5971 2202
rect 6023 2150 6035 2202
rect 6087 2150 8194 2202
rect 8246 2150 8258 2202
rect 8310 2150 8322 2202
rect 8374 2150 8386 2202
rect 8438 2150 8450 2202
rect 8502 2150 10609 2202
rect 10661 2150 10673 2202
rect 10725 2150 10737 2202
rect 10789 2150 10801 2202
rect 10853 2150 10865 2202
rect 10917 2150 10923 2202
rect 1104 2128 10923 2150
<< via1 >>
rect 2157 11398 2209 11450
rect 2221 11398 2273 11450
rect 2285 11398 2337 11450
rect 2349 11398 2401 11450
rect 2413 11398 2465 11450
rect 4572 11398 4624 11450
rect 4636 11398 4688 11450
rect 4700 11398 4752 11450
rect 4764 11398 4816 11450
rect 4828 11398 4880 11450
rect 6987 11398 7039 11450
rect 7051 11398 7103 11450
rect 7115 11398 7167 11450
rect 7179 11398 7231 11450
rect 7243 11398 7295 11450
rect 9402 11398 9454 11450
rect 9466 11398 9518 11450
rect 9530 11398 9582 11450
rect 9594 11398 9646 11450
rect 9658 11398 9710 11450
rect 2964 11296 3016 11348
rect 8944 11296 8996 11348
rect 4252 11092 4304 11144
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 3148 11024 3200 11033
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 7380 11024 7432 11076
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 3240 10956 3292 11008
rect 7932 10956 7984 11008
rect 3364 10854 3416 10906
rect 3428 10854 3480 10906
rect 3492 10854 3544 10906
rect 3556 10854 3608 10906
rect 3620 10854 3672 10906
rect 5779 10854 5831 10906
rect 5843 10854 5895 10906
rect 5907 10854 5959 10906
rect 5971 10854 6023 10906
rect 6035 10854 6087 10906
rect 8194 10854 8246 10906
rect 8258 10854 8310 10906
rect 8322 10854 8374 10906
rect 8386 10854 8438 10906
rect 8450 10854 8502 10906
rect 10609 10854 10661 10906
rect 10673 10854 10725 10906
rect 10737 10854 10789 10906
rect 10801 10854 10853 10906
rect 10865 10854 10917 10906
rect 3148 10752 3200 10804
rect 940 10616 992 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 8116 10752 8168 10804
rect 9128 10752 9180 10804
rect 8392 10684 8444 10736
rect 4436 10548 4488 10600
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 6920 10616 6972 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7748 10616 7800 10668
rect 8852 10616 8904 10668
rect 7840 10548 7892 10600
rect 10876 10480 10928 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 3884 10412 3936 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5724 10412 5776 10464
rect 6828 10412 6880 10464
rect 6920 10412 6972 10464
rect 7564 10412 7616 10464
rect 7656 10412 7708 10464
rect 9220 10412 9272 10464
rect 2157 10310 2209 10362
rect 2221 10310 2273 10362
rect 2285 10310 2337 10362
rect 2349 10310 2401 10362
rect 2413 10310 2465 10362
rect 4572 10310 4624 10362
rect 4636 10310 4688 10362
rect 4700 10310 4752 10362
rect 4764 10310 4816 10362
rect 4828 10310 4880 10362
rect 6987 10310 7039 10362
rect 7051 10310 7103 10362
rect 7115 10310 7167 10362
rect 7179 10310 7231 10362
rect 7243 10310 7295 10362
rect 9402 10310 9454 10362
rect 9466 10310 9518 10362
rect 9530 10310 9582 10362
rect 9594 10310 9646 10362
rect 9658 10310 9710 10362
rect 1584 10208 1636 10260
rect 3240 10251 3292 10260
rect 3240 10217 3249 10251
rect 3249 10217 3283 10251
rect 3283 10217 3292 10251
rect 3240 10208 3292 10217
rect 3424 10208 3476 10260
rect 5540 10208 5592 10260
rect 5724 10208 5776 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 7380 10140 7432 10192
rect 3700 10004 3752 10056
rect 5632 10004 5684 10056
rect 3884 9936 3936 9988
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 8208 10208 8260 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 7932 10140 7984 10192
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 3792 9868 3844 9920
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 6552 9979 6604 9988
rect 6552 9945 6586 9979
rect 6586 9945 6604 9979
rect 6552 9936 6604 9945
rect 7656 9936 7708 9988
rect 6000 9868 6052 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8668 10072 8720 10124
rect 9220 10072 9272 10124
rect 10416 10208 10468 10260
rect 9496 9868 9548 9920
rect 3364 9766 3416 9818
rect 3428 9766 3480 9818
rect 3492 9766 3544 9818
rect 3556 9766 3608 9818
rect 3620 9766 3672 9818
rect 5779 9766 5831 9818
rect 5843 9766 5895 9818
rect 5907 9766 5959 9818
rect 5971 9766 6023 9818
rect 6035 9766 6087 9818
rect 8194 9766 8246 9818
rect 8258 9766 8310 9818
rect 8322 9766 8374 9818
rect 8386 9766 8438 9818
rect 8450 9766 8502 9818
rect 10609 9766 10661 9818
rect 10673 9766 10725 9818
rect 10737 9766 10789 9818
rect 10801 9766 10853 9818
rect 10865 9766 10917 9818
rect 3700 9528 3752 9580
rect 5172 9664 5224 9716
rect 5264 9664 5316 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7472 9528 7524 9580
rect 7748 9528 7800 9580
rect 8668 9664 8720 9716
rect 9496 9596 9548 9648
rect 4436 9460 4488 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 6828 9460 6880 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 4252 9392 4304 9444
rect 5448 9392 5500 9444
rect 6000 9324 6052 9376
rect 7380 9324 7432 9376
rect 7932 9324 7984 9376
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 2157 9222 2209 9274
rect 2221 9222 2273 9274
rect 2285 9222 2337 9274
rect 2349 9222 2401 9274
rect 2413 9222 2465 9274
rect 4572 9222 4624 9274
rect 4636 9222 4688 9274
rect 4700 9222 4752 9274
rect 4764 9222 4816 9274
rect 4828 9222 4880 9274
rect 6987 9222 7039 9274
rect 7051 9222 7103 9274
rect 7115 9222 7167 9274
rect 7179 9222 7231 9274
rect 7243 9222 7295 9274
rect 9402 9222 9454 9274
rect 9466 9222 9518 9274
rect 9530 9222 9582 9274
rect 9594 9222 9646 9274
rect 9658 9222 9710 9274
rect 3608 9120 3660 9172
rect 4436 9120 4488 9172
rect 5080 9120 5132 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 5448 8984 5500 9036
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6736 9052 6788 9104
rect 7840 9052 7892 9104
rect 5632 8848 5684 8900
rect 7288 8848 7340 8900
rect 7564 8848 7616 8900
rect 7748 8848 7800 8900
rect 7932 8848 7984 8900
rect 8024 8891 8076 8900
rect 8024 8857 8033 8891
rect 8033 8857 8067 8891
rect 8067 8857 8076 8891
rect 8024 8848 8076 8857
rect 9864 8848 9916 8900
rect 9220 8780 9272 8832
rect 3364 8678 3416 8730
rect 3428 8678 3480 8730
rect 3492 8678 3544 8730
rect 3556 8678 3608 8730
rect 3620 8678 3672 8730
rect 5779 8678 5831 8730
rect 5843 8678 5895 8730
rect 5907 8678 5959 8730
rect 5971 8678 6023 8730
rect 6035 8678 6087 8730
rect 8194 8678 8246 8730
rect 8258 8678 8310 8730
rect 8322 8678 8374 8730
rect 8386 8678 8438 8730
rect 8450 8678 8502 8730
rect 10609 8678 10661 8730
rect 10673 8678 10725 8730
rect 10737 8678 10789 8730
rect 10801 8678 10853 8730
rect 10865 8678 10917 8730
rect 7656 8576 7708 8628
rect 8024 8576 8076 8628
rect 8116 8576 8168 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 3700 8440 3752 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 6368 8372 6420 8424
rect 6828 8372 6880 8424
rect 3976 8304 4028 8356
rect 7840 8304 7892 8356
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 5540 8236 5592 8288
rect 6828 8236 6880 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 2157 8134 2209 8186
rect 2221 8134 2273 8186
rect 2285 8134 2337 8186
rect 2349 8134 2401 8186
rect 2413 8134 2465 8186
rect 4572 8134 4624 8186
rect 4636 8134 4688 8186
rect 4700 8134 4752 8186
rect 4764 8134 4816 8186
rect 4828 8134 4880 8186
rect 6987 8134 7039 8186
rect 7051 8134 7103 8186
rect 7115 8134 7167 8186
rect 7179 8134 7231 8186
rect 7243 8134 7295 8186
rect 9402 8134 9454 8186
rect 9466 8134 9518 8186
rect 9530 8134 9582 8186
rect 9594 8134 9646 8186
rect 9658 8134 9710 8186
rect 1860 8032 1912 8084
rect 7472 8032 7524 8084
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 6828 7964 6880 8016
rect 9128 7964 9180 8016
rect 2872 7896 2924 7948
rect 2964 7896 3016 7948
rect 3884 7896 3936 7948
rect 3240 7760 3292 7812
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 6184 7760 6236 7812
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 3792 7692 3844 7744
rect 6368 7692 6420 7744
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9772 7692 9824 7744
rect 9956 7692 10008 7744
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 10232 7692 10284 7744
rect 10324 7692 10376 7744
rect 3364 7590 3416 7642
rect 3428 7590 3480 7642
rect 3492 7590 3544 7642
rect 3556 7590 3608 7642
rect 3620 7590 3672 7642
rect 5779 7590 5831 7642
rect 5843 7590 5895 7642
rect 5907 7590 5959 7642
rect 5971 7590 6023 7642
rect 6035 7590 6087 7642
rect 8194 7590 8246 7642
rect 8258 7590 8310 7642
rect 8322 7590 8374 7642
rect 8386 7590 8438 7642
rect 8450 7590 8502 7642
rect 10609 7590 10661 7642
rect 10673 7590 10725 7642
rect 10737 7590 10789 7642
rect 10801 7590 10853 7642
rect 10865 7590 10917 7642
rect 1584 7488 1636 7540
rect 3608 7352 3660 7404
rect 3792 7488 3844 7540
rect 5540 7420 5592 7472
rect 7472 7488 7524 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 8576 7488 8628 7540
rect 8944 7488 8996 7540
rect 9128 7488 9180 7540
rect 9220 7488 9272 7540
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2964 7284 3016 7336
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 3608 7148 3660 7200
rect 5632 7352 5684 7404
rect 8024 7420 8076 7472
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 7840 7284 7892 7336
rect 8576 7284 8628 7336
rect 8668 7216 8720 7268
rect 10324 7463 10376 7472
rect 10324 7429 10333 7463
rect 10333 7429 10367 7463
rect 10367 7429 10376 7463
rect 10324 7420 10376 7429
rect 9312 7352 9364 7404
rect 10232 7352 10284 7404
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 2157 7046 2209 7098
rect 2221 7046 2273 7098
rect 2285 7046 2337 7098
rect 2349 7046 2401 7098
rect 2413 7046 2465 7098
rect 4572 7046 4624 7098
rect 4636 7046 4688 7098
rect 4700 7046 4752 7098
rect 4764 7046 4816 7098
rect 4828 7046 4880 7098
rect 6987 7046 7039 7098
rect 7051 7046 7103 7098
rect 7115 7046 7167 7098
rect 7179 7046 7231 7098
rect 7243 7046 7295 7098
rect 9402 7046 9454 7098
rect 9466 7046 9518 7098
rect 9530 7046 9582 7098
rect 9594 7046 9646 7098
rect 9658 7046 9710 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 2872 6944 2924 6996
rect 3884 6944 3936 6996
rect 8576 6944 8628 6996
rect 9312 6876 9364 6928
rect 1860 6808 1912 6860
rect 5540 6808 5592 6860
rect 9864 6808 9916 6860
rect 2964 6740 3016 6792
rect 3240 6740 3292 6792
rect 3424 6672 3476 6724
rect 4160 6672 4212 6724
rect 7748 6672 7800 6724
rect 2780 6604 2832 6656
rect 6184 6604 6236 6656
rect 8576 6604 8628 6656
rect 8852 6604 8904 6656
rect 3364 6502 3416 6554
rect 3428 6502 3480 6554
rect 3492 6502 3544 6554
rect 3556 6502 3608 6554
rect 3620 6502 3672 6554
rect 5779 6502 5831 6554
rect 5843 6502 5895 6554
rect 5907 6502 5959 6554
rect 5971 6502 6023 6554
rect 6035 6502 6087 6554
rect 8194 6502 8246 6554
rect 8258 6502 8310 6554
rect 8322 6502 8374 6554
rect 8386 6502 8438 6554
rect 8450 6502 8502 6554
rect 10609 6502 10661 6554
rect 10673 6502 10725 6554
rect 10737 6502 10789 6554
rect 10801 6502 10853 6554
rect 10865 6502 10917 6554
rect 7748 6443 7800 6452
rect 7748 6409 7757 6443
rect 7757 6409 7791 6443
rect 7791 6409 7800 6443
rect 7748 6400 7800 6409
rect 7932 6400 7984 6452
rect 8852 6400 8904 6452
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 5264 6264 5316 6316
rect 5632 6264 5684 6316
rect 10232 6400 10284 6452
rect 3240 6196 3292 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 8668 6264 8720 6316
rect 5540 6060 5592 6112
rect 5816 6060 5868 6112
rect 6276 6060 6328 6112
rect 8576 6060 8628 6112
rect 2157 5958 2209 6010
rect 2221 5958 2273 6010
rect 2285 5958 2337 6010
rect 2349 5958 2401 6010
rect 2413 5958 2465 6010
rect 4572 5958 4624 6010
rect 4636 5958 4688 6010
rect 4700 5958 4752 6010
rect 4764 5958 4816 6010
rect 4828 5958 4880 6010
rect 6987 5958 7039 6010
rect 7051 5958 7103 6010
rect 7115 5958 7167 6010
rect 7179 5958 7231 6010
rect 7243 5958 7295 6010
rect 9402 5958 9454 6010
rect 9466 5958 9518 6010
rect 9530 5958 9582 6010
rect 9594 5958 9646 6010
rect 9658 5958 9710 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 3240 5856 3292 5908
rect 7656 5856 7708 5908
rect 8852 5856 8904 5908
rect 9772 5856 9824 5908
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 2780 5695 2832 5704
rect 2780 5661 2789 5695
rect 2789 5661 2823 5695
rect 2823 5661 2832 5695
rect 2780 5652 2832 5661
rect 3976 5652 4028 5704
rect 6276 5584 6328 5636
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 2228 5516 2280 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 5264 5559 5316 5568
rect 5264 5525 5273 5559
rect 5273 5525 5307 5559
rect 5307 5525 5316 5559
rect 5264 5516 5316 5525
rect 5632 5516 5684 5568
rect 7840 5516 7892 5568
rect 9036 5516 9088 5568
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 3364 5414 3416 5466
rect 3428 5414 3480 5466
rect 3492 5414 3544 5466
rect 3556 5414 3608 5466
rect 3620 5414 3672 5466
rect 5779 5414 5831 5466
rect 5843 5414 5895 5466
rect 5907 5414 5959 5466
rect 5971 5414 6023 5466
rect 6035 5414 6087 5466
rect 8194 5414 8246 5466
rect 8258 5414 8310 5466
rect 8322 5414 8374 5466
rect 8386 5414 8438 5466
rect 8450 5414 8502 5466
rect 10609 5414 10661 5466
rect 10673 5414 10725 5466
rect 10737 5414 10789 5466
rect 10801 5414 10853 5466
rect 10865 5414 10917 5466
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 4712 5312 4764 5364
rect 6276 5312 6328 5364
rect 5540 5244 5592 5296
rect 9220 5244 9272 5296
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 2688 5108 2740 5160
rect 3240 5108 3292 5160
rect 8576 5176 8628 5228
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 5632 4972 5684 5024
rect 8760 4972 8812 5024
rect 9128 4972 9180 5024
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 2157 4870 2209 4922
rect 2221 4870 2273 4922
rect 2285 4870 2337 4922
rect 2349 4870 2401 4922
rect 2413 4870 2465 4922
rect 4572 4870 4624 4922
rect 4636 4870 4688 4922
rect 4700 4870 4752 4922
rect 4764 4870 4816 4922
rect 4828 4870 4880 4922
rect 6987 4870 7039 4922
rect 7051 4870 7103 4922
rect 7115 4870 7167 4922
rect 7179 4870 7231 4922
rect 7243 4870 7295 4922
rect 9402 4870 9454 4922
rect 9466 4870 9518 4922
rect 9530 4870 9582 4922
rect 9594 4870 9646 4922
rect 9658 4870 9710 4922
rect 3700 4768 3752 4820
rect 7564 4700 7616 4752
rect 9772 4768 9824 4820
rect 8852 4700 8904 4752
rect 8668 4675 8720 4684
rect 8668 4641 8677 4675
rect 8677 4641 8711 4675
rect 8711 4641 8720 4675
rect 8668 4632 8720 4641
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 9864 4632 9916 4684
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 9036 4564 9088 4616
rect 9220 4564 9272 4616
rect 4436 4428 4488 4480
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 3364 4326 3416 4378
rect 3428 4326 3480 4378
rect 3492 4326 3544 4378
rect 3556 4326 3608 4378
rect 3620 4326 3672 4378
rect 5779 4326 5831 4378
rect 5843 4326 5895 4378
rect 5907 4326 5959 4378
rect 5971 4326 6023 4378
rect 6035 4326 6087 4378
rect 8194 4326 8246 4378
rect 8258 4326 8310 4378
rect 8322 4326 8374 4378
rect 8386 4326 8438 4378
rect 8450 4326 8502 4378
rect 10609 4326 10661 4378
rect 10673 4326 10725 4378
rect 10737 4326 10789 4378
rect 10801 4326 10853 4378
rect 10865 4326 10917 4378
rect 7288 4224 7340 4276
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3976 4020 4028 4072
rect 5540 4088 5592 4140
rect 4436 4020 4488 4072
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 7748 4088 7800 4140
rect 8024 4088 8076 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9864 4088 9916 4140
rect 10048 4088 10100 4140
rect 2688 3884 2740 3936
rect 5264 3952 5316 4004
rect 8208 3952 8260 4004
rect 5724 3884 5776 3936
rect 8852 4020 8904 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 9220 3884 9272 3936
rect 2157 3782 2209 3834
rect 2221 3782 2273 3834
rect 2285 3782 2337 3834
rect 2349 3782 2401 3834
rect 2413 3782 2465 3834
rect 4572 3782 4624 3834
rect 4636 3782 4688 3834
rect 4700 3782 4752 3834
rect 4764 3782 4816 3834
rect 4828 3782 4880 3834
rect 6987 3782 7039 3834
rect 7051 3782 7103 3834
rect 7115 3782 7167 3834
rect 7179 3782 7231 3834
rect 7243 3782 7295 3834
rect 9402 3782 9454 3834
rect 9466 3782 9518 3834
rect 9530 3782 9582 3834
rect 9594 3782 9646 3834
rect 9658 3782 9710 3834
rect 3332 3680 3384 3732
rect 5724 3680 5776 3732
rect 7748 3680 7800 3732
rect 8668 3680 8720 3732
rect 9956 3680 10008 3732
rect 10324 3680 10376 3732
rect 1952 3544 2004 3596
rect 5632 3544 5684 3596
rect 3240 3476 3292 3528
rect 3700 3476 3752 3528
rect 8576 3544 8628 3596
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 5448 3408 5500 3460
rect 5540 3340 5592 3392
rect 6276 3340 6328 3392
rect 8208 3476 8260 3528
rect 7932 3408 7984 3460
rect 7288 3340 7340 3392
rect 7748 3340 7800 3392
rect 9128 3476 9180 3528
rect 9864 3408 9916 3460
rect 3364 3238 3416 3290
rect 3428 3238 3480 3290
rect 3492 3238 3544 3290
rect 3556 3238 3608 3290
rect 3620 3238 3672 3290
rect 5779 3238 5831 3290
rect 5843 3238 5895 3290
rect 5907 3238 5959 3290
rect 5971 3238 6023 3290
rect 6035 3238 6087 3290
rect 8194 3238 8246 3290
rect 8258 3238 8310 3290
rect 8322 3238 8374 3290
rect 8386 3238 8438 3290
rect 8450 3238 8502 3290
rect 10609 3238 10661 3290
rect 10673 3238 10725 3290
rect 10737 3238 10789 3290
rect 10801 3238 10853 3290
rect 10865 3238 10917 3290
rect 1860 3136 1912 3188
rect 3792 3136 3844 3188
rect 2872 3000 2924 3052
rect 6184 3111 6236 3120
rect 6184 3077 6193 3111
rect 6193 3077 6227 3111
rect 6227 3077 6236 3111
rect 6184 3068 6236 3077
rect 7840 3136 7892 3188
rect 8392 3136 8444 3188
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10416 3136 10468 3188
rect 7288 3068 7340 3120
rect 5540 2932 5592 2984
rect 3240 2864 3292 2916
rect 4068 2864 4120 2916
rect 3700 2796 3752 2848
rect 7748 3000 7800 3052
rect 7932 3043 7984 3052
rect 7932 3009 7966 3043
rect 7966 3009 7984 3043
rect 7932 3000 7984 3009
rect 10876 3000 10928 3052
rect 7564 2864 7616 2916
rect 9772 2796 9824 2848
rect 2157 2694 2209 2746
rect 2221 2694 2273 2746
rect 2285 2694 2337 2746
rect 2349 2694 2401 2746
rect 2413 2694 2465 2746
rect 4572 2694 4624 2746
rect 4636 2694 4688 2746
rect 4700 2694 4752 2746
rect 4764 2694 4816 2746
rect 4828 2694 4880 2746
rect 6987 2694 7039 2746
rect 7051 2694 7103 2746
rect 7115 2694 7167 2746
rect 7179 2694 7231 2746
rect 7243 2694 7295 2746
rect 9402 2694 9454 2746
rect 9466 2694 9518 2746
rect 9530 2694 9582 2746
rect 9594 2694 9646 2746
rect 9658 2694 9710 2746
rect 2872 2592 2924 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 7564 2592 7616 2644
rect 7932 2592 7984 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 8392 2567 8444 2576
rect 8392 2533 8401 2567
rect 8401 2533 8435 2567
rect 8435 2533 8444 2567
rect 8392 2524 8444 2533
rect 3700 2456 3752 2508
rect 9036 2456 9088 2508
rect 10324 2499 10376 2508
rect 10324 2465 10333 2499
rect 10333 2465 10367 2499
rect 10367 2465 10376 2499
rect 10324 2456 10376 2465
rect 2964 2388 3016 2440
rect 3976 2320 4028 2372
rect 4160 2320 4212 2372
rect 8116 2388 8168 2440
rect 8760 2320 8812 2372
rect 5448 2252 5500 2304
rect 8944 2252 8996 2304
rect 3364 2150 3416 2202
rect 3428 2150 3480 2202
rect 3492 2150 3544 2202
rect 3556 2150 3608 2202
rect 3620 2150 3672 2202
rect 5779 2150 5831 2202
rect 5843 2150 5895 2202
rect 5907 2150 5959 2202
rect 5971 2150 6023 2202
rect 6035 2150 6087 2202
rect 8194 2150 8246 2202
rect 8258 2150 8310 2202
rect 8322 2150 8374 2202
rect 8386 2150 8438 2202
rect 8450 2150 8502 2202
rect 10609 2150 10661 2202
rect 10673 2150 10725 2202
rect 10737 2150 10789 2202
rect 10801 2150 10853 2202
rect 10865 2150 10917 2202
<< metal2 >>
rect 2962 13298 3018 14098
rect 8942 13298 8998 14098
rect 2157 11452 2465 11461
rect 2157 11450 2163 11452
rect 2219 11450 2243 11452
rect 2299 11450 2323 11452
rect 2379 11450 2403 11452
rect 2459 11450 2465 11452
rect 2219 11398 2221 11450
rect 2401 11398 2403 11450
rect 2157 11396 2163 11398
rect 2219 11396 2243 11398
rect 2299 11396 2323 11398
rect 2379 11396 2403 11398
rect 2459 11396 2465 11398
rect 2157 11387 2465 11396
rect 2976 11354 3004 13298
rect 4572 11452 4880 11461
rect 4572 11450 4578 11452
rect 4634 11450 4658 11452
rect 4714 11450 4738 11452
rect 4794 11450 4818 11452
rect 4874 11450 4880 11452
rect 4634 11398 4636 11450
rect 4816 11398 4818 11450
rect 4572 11396 4578 11398
rect 4634 11396 4658 11398
rect 4714 11396 4738 11398
rect 4794 11396 4818 11398
rect 4874 11396 4880 11398
rect 4572 11387 4880 11396
rect 6987 11452 7295 11461
rect 6987 11450 6993 11452
rect 7049 11450 7073 11452
rect 7129 11450 7153 11452
rect 7209 11450 7233 11452
rect 7289 11450 7295 11452
rect 7049 11398 7051 11450
rect 7231 11398 7233 11450
rect 6987 11396 6993 11398
rect 7049 11396 7073 11398
rect 7129 11396 7153 11398
rect 7209 11396 7233 11398
rect 7289 11396 7295 11398
rect 6987 11387 7295 11396
rect 8956 11354 8984 13298
rect 9402 11452 9710 11461
rect 9402 11450 9408 11452
rect 9464 11450 9488 11452
rect 9544 11450 9568 11452
rect 9624 11450 9648 11452
rect 9704 11450 9710 11452
rect 9464 11398 9466 11450
rect 9646 11398 9648 11450
rect 9402 11396 9408 11398
rect 9464 11396 9488 11398
rect 9544 11396 9568 11398
rect 9624 11396 9648 11398
rect 9704 11396 9710 11398
rect 9402 11387 9710 11396
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3160 10810 3188 11018
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 952 10441 980 10610
rect 1584 10464 1636 10470
rect 938 10432 994 10441
rect 1584 10406 1636 10412
rect 938 10367 994 10376
rect 1596 10266 1624 10406
rect 2157 10364 2465 10373
rect 2157 10362 2163 10364
rect 2219 10362 2243 10364
rect 2299 10362 2323 10364
rect 2379 10362 2403 10364
rect 2459 10362 2465 10364
rect 2219 10310 2221 10362
rect 2401 10310 2403 10362
rect 2157 10308 2163 10310
rect 2219 10308 2243 10310
rect 2299 10308 2323 10310
rect 2379 10308 2403 10310
rect 2459 10308 2465 10310
rect 2157 10299 2465 10308
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 2157 9276 2465 9285
rect 2157 9274 2163 9276
rect 2219 9274 2243 9276
rect 2299 9274 2323 9276
rect 2379 9274 2403 9276
rect 2459 9274 2465 9276
rect 2219 9222 2221 9274
rect 2401 9222 2403 9274
rect 2157 9220 2163 9222
rect 2219 9220 2243 9222
rect 2299 9220 2323 9222
rect 2379 9220 2403 9222
rect 2459 9220 2465 9222
rect 2157 9211 2465 9220
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 7546 1624 8434
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 8090 1900 8366
rect 2157 8188 2465 8197
rect 2157 8186 2163 8188
rect 2219 8186 2243 8188
rect 2299 8186 2323 8188
rect 2379 8186 2403 8188
rect 2459 8186 2465 8188
rect 2219 8134 2221 8186
rect 2401 8134 2403 8186
rect 2157 8132 2163 8134
rect 2219 8132 2243 8134
rect 2299 8132 2323 8134
rect 2379 8132 2403 8134
rect 2459 8132 2465 8134
rect 2157 8123 2465 8132
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 7002 1992 7278
rect 2157 7100 2465 7109
rect 2157 7098 2163 7100
rect 2219 7098 2243 7100
rect 2299 7098 2323 7100
rect 2379 7098 2403 7100
rect 2459 7098 2465 7100
rect 2219 7046 2221 7098
rect 2401 7046 2403 7098
rect 2157 7044 2163 7046
rect 2219 7044 2243 7046
rect 2299 7044 2323 7046
rect 2379 7044 2403 7046
rect 2459 7044 2465 7046
rect 2157 7035 2465 7044
rect 2884 7002 2912 7890
rect 2976 7342 3004 7890
rect 3068 7562 3096 10610
rect 3252 10266 3280 10950
rect 3364 10908 3672 10917
rect 3364 10906 3370 10908
rect 3426 10906 3450 10908
rect 3506 10906 3530 10908
rect 3586 10906 3610 10908
rect 3666 10906 3672 10908
rect 3426 10854 3428 10906
rect 3608 10854 3610 10906
rect 3364 10852 3370 10854
rect 3426 10852 3450 10854
rect 3506 10852 3530 10854
rect 3586 10852 3610 10854
rect 3666 10852 3672 10854
rect 3364 10843 3672 10852
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 10266 3464 10610
rect 4264 10470 4292 11086
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 5779 10908 6087 10917
rect 5779 10906 5785 10908
rect 5841 10906 5865 10908
rect 5921 10906 5945 10908
rect 6001 10906 6025 10908
rect 6081 10906 6087 10908
rect 5841 10854 5843 10906
rect 6023 10854 6025 10906
rect 5779 10852 5785 10854
rect 5841 10852 5865 10854
rect 5921 10852 5945 10854
rect 6001 10852 6025 10854
rect 6081 10852 6087 10854
rect 5779 10843 6087 10852
rect 6932 10674 6960 11018
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3364 9820 3672 9829
rect 3364 9818 3370 9820
rect 3426 9818 3450 9820
rect 3506 9818 3530 9820
rect 3586 9818 3610 9820
rect 3666 9818 3672 9820
rect 3426 9766 3428 9818
rect 3608 9766 3610 9818
rect 3364 9764 3370 9766
rect 3426 9764 3450 9766
rect 3506 9764 3530 9766
rect 3586 9764 3610 9766
rect 3666 9764 3672 9766
rect 3364 9755 3672 9764
rect 3712 9586 3740 9998
rect 3896 9994 3924 10406
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9178 3648 9318
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3364 8732 3672 8741
rect 3364 8730 3370 8732
rect 3426 8730 3450 8732
rect 3506 8730 3530 8732
rect 3586 8730 3610 8732
rect 3666 8730 3672 8732
rect 3426 8678 3428 8730
rect 3608 8678 3610 8730
rect 3364 8676 3370 8678
rect 3426 8676 3450 8678
rect 3506 8676 3530 8678
rect 3586 8676 3610 8678
rect 3666 8676 3672 8678
rect 3364 8667 3672 8676
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3068 7534 3188 7562
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 5914 1900 6802
rect 2976 6798 3004 7278
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2157 6012 2465 6021
rect 2157 6010 2163 6012
rect 2219 6010 2243 6012
rect 2299 6010 2323 6012
rect 2379 6010 2403 6012
rect 2459 6010 2465 6012
rect 2219 5958 2221 6010
rect 2401 5958 2403 6010
rect 2157 5956 2163 5958
rect 2219 5956 2243 5958
rect 2299 5956 2323 5958
rect 2379 5956 2403 5958
rect 2459 5956 2465 5958
rect 2157 5947 2465 5956
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2792 5710 2820 6598
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 5166 2268 5510
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1964 3602 1992 5102
rect 2157 4924 2465 4933
rect 2157 4922 2163 4924
rect 2219 4922 2243 4924
rect 2299 4922 2323 4924
rect 2379 4922 2403 4924
rect 2459 4922 2465 4924
rect 2219 4870 2221 4922
rect 2401 4870 2403 4922
rect 2157 4868 2163 4870
rect 2219 4868 2243 4870
rect 2299 4868 2323 4870
rect 2379 4868 2403 4870
rect 2459 4868 2465 4870
rect 2157 4859 2465 4868
rect 2700 3942 2728 5102
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2157 3836 2465 3845
rect 2157 3834 2163 3836
rect 2219 3834 2243 3836
rect 2299 3834 2323 3836
rect 2379 3834 2403 3836
rect 2459 3834 2465 3836
rect 2219 3782 2221 3834
rect 2401 3782 2403 3834
rect 2157 3780 2163 3782
rect 2219 3780 2243 3782
rect 2299 3780 2323 3782
rect 2379 3780 2403 3782
rect 2459 3780 2465 3782
rect 2157 3771 2465 3780
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1872 3194 1900 3402
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2884 3058 2912 5714
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3160 2774 3188 7534
rect 3252 6798 3280 7754
rect 3364 7644 3672 7653
rect 3364 7642 3370 7644
rect 3426 7642 3450 7644
rect 3506 7642 3530 7644
rect 3586 7642 3610 7644
rect 3666 7642 3672 7644
rect 3426 7590 3428 7642
rect 3608 7590 3610 7642
rect 3364 7588 3370 7590
rect 3426 7588 3450 7590
rect 3506 7588 3530 7590
rect 3586 7588 3610 7590
rect 3666 7588 3672 7590
rect 3364 7579 3672 7588
rect 3712 7426 3740 8434
rect 3804 7750 3832 9862
rect 4264 9450 4292 10406
rect 4448 9518 4476 10542
rect 4572 10364 4880 10373
rect 4572 10362 4578 10364
rect 4634 10362 4658 10364
rect 4714 10362 4738 10364
rect 4794 10362 4818 10364
rect 4874 10362 4880 10364
rect 4634 10310 4636 10362
rect 4816 10310 4818 10362
rect 4572 10308 4578 10310
rect 4634 10308 4658 10310
rect 4714 10308 4738 10310
rect 4794 10308 4818 10310
rect 4874 10308 4880 10310
rect 4572 10299 4880 10308
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5184 9722 5212 9862
rect 5276 9722 5304 9862
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4448 9178 4476 9454
rect 4572 9276 4880 9285
rect 4572 9274 4578 9276
rect 4634 9274 4658 9276
rect 4714 9274 4738 9276
rect 4794 9274 4818 9276
rect 4874 9274 4880 9276
rect 4634 9222 4636 9274
rect 4816 9222 4818 9274
rect 4572 9220 4578 9222
rect 4634 9220 4658 9222
rect 4714 9220 4738 9222
rect 4794 9220 4818 9222
rect 4874 9220 4880 9222
rect 4572 9211 4880 9220
rect 5092 9178 5120 9454
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5460 9042 5488 9386
rect 5552 9178 5580 10202
rect 5644 10062 5672 10542
rect 6932 10470 6960 10610
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 5736 10266 5764 10406
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9926 6040 9998
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5779 9820 6087 9829
rect 5779 9818 5785 9820
rect 5841 9818 5865 9820
rect 5921 9818 5945 9820
rect 6001 9818 6025 9820
rect 6081 9818 6087 9820
rect 5841 9766 5843 9818
rect 6023 9766 6025 9818
rect 5779 9764 5785 9766
rect 5841 9764 5865 9766
rect 5921 9764 5945 9766
rect 6001 9764 6025 9766
rect 6081 9764 6087 9766
rect 5779 9755 6087 9764
rect 6564 9722 6592 9930
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 6012 8974 6040 9318
rect 6748 9110 6776 9658
rect 6840 9602 6868 10406
rect 6987 10364 7295 10373
rect 6987 10362 6993 10364
rect 7049 10362 7073 10364
rect 7129 10362 7153 10364
rect 7209 10362 7233 10364
rect 7289 10362 7295 10364
rect 7049 10310 7051 10362
rect 7231 10310 7233 10362
rect 6987 10308 6993 10310
rect 7049 10308 7073 10310
rect 7129 10308 7153 10310
rect 7209 10308 7233 10310
rect 7289 10308 7295 10310
rect 6987 10299 7295 10308
rect 7392 10198 7420 11018
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 6840 9586 7328 9602
rect 7392 9586 7420 10134
rect 7484 9586 7512 10610
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7576 9722 7604 10406
rect 7668 10266 7696 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7760 10010 7788 10610
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7668 9994 7788 10010
rect 7656 9988 7788 9994
rect 7708 9982 7788 9988
rect 7656 9930 7708 9936
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 6840 9580 7340 9586
rect 6840 9574 7288 9580
rect 7288 9522 7340 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 7104 9512 7156 9518
rect 7156 9460 7420 9466
rect 7104 9454 7420 9460
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7954 3924 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7546 3832 7686
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3620 7410 3740 7426
rect 3608 7404 3740 7410
rect 3660 7398 3740 7404
rect 3608 7346 3660 7352
rect 3620 7206 3648 7346
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6254 3280 6734
rect 3436 6730 3464 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3364 6556 3672 6565
rect 3364 6554 3370 6556
rect 3426 6554 3450 6556
rect 3506 6554 3530 6556
rect 3586 6554 3610 6556
rect 3666 6554 3672 6556
rect 3426 6502 3428 6554
rect 3608 6502 3610 6554
rect 3364 6500 3370 6502
rect 3426 6500 3450 6502
rect 3506 6500 3530 6502
rect 3586 6500 3610 6502
rect 3666 6500 3672 6502
rect 3364 6491 3672 6500
rect 3896 6254 3924 6938
rect 3988 6322 4016 8298
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 4572 8188 4880 8197
rect 4572 8186 4578 8188
rect 4634 8186 4658 8188
rect 4714 8186 4738 8188
rect 4794 8186 4818 8188
rect 4874 8186 4880 8188
rect 4634 8134 4636 8186
rect 4816 8134 4818 8186
rect 4572 8132 4578 8134
rect 4634 8132 4658 8134
rect 4714 8132 4738 8134
rect 4794 8132 4818 8134
rect 4874 8132 4880 8134
rect 4572 8123 4880 8132
rect 5552 7478 5580 8230
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5644 7410 5672 8842
rect 5779 8732 6087 8741
rect 5779 8730 5785 8732
rect 5841 8730 5865 8732
rect 5921 8730 5945 8732
rect 6001 8730 6025 8732
rect 6081 8730 6087 8732
rect 5841 8678 5843 8730
rect 6023 8678 6025 8730
rect 5779 8676 5785 8678
rect 5841 8676 5865 8678
rect 5921 8676 5945 8678
rect 6001 8676 6025 8678
rect 6081 8676 6087 8678
rect 5779 8667 6087 8676
rect 6840 8430 6868 9454
rect 7116 9438 7420 9454
rect 7392 9382 7420 9438
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 6987 9276 7295 9285
rect 6987 9274 6993 9276
rect 7049 9274 7073 9276
rect 7129 9274 7153 9276
rect 7209 9274 7233 9276
rect 7289 9274 7295 9276
rect 7049 9222 7051 9274
rect 7231 9222 7233 9274
rect 6987 9220 6993 9222
rect 7049 9220 7073 9222
rect 7129 9220 7153 9222
rect 7209 9220 7233 9222
rect 7289 9220 7295 9222
rect 6987 9211 7295 9220
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8498 7328 8842
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 5779 7644 6087 7653
rect 5779 7642 5785 7644
rect 5841 7642 5865 7644
rect 5921 7642 5945 7644
rect 6001 7642 6025 7644
rect 6081 7642 6087 7644
rect 5841 7590 5843 7642
rect 6023 7590 6025 7642
rect 5779 7588 5785 7590
rect 5841 7588 5865 7590
rect 5921 7588 5945 7590
rect 6001 7588 6025 7590
rect 6081 7588 6087 7590
rect 5779 7579 6087 7588
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 4572 7100 4880 7109
rect 4572 7098 4578 7100
rect 4634 7098 4658 7100
rect 4714 7098 4738 7100
rect 4794 7098 4818 7100
rect 4874 7098 4880 7100
rect 4634 7046 4636 7098
rect 4816 7046 4818 7098
rect 4572 7044 4578 7046
rect 4634 7044 4658 7046
rect 4714 7044 4738 7046
rect 4794 7044 4818 7046
rect 4874 7044 4880 7046
rect 4572 7035 4880 7044
rect 5552 6866 5580 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3252 5914 3280 6190
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3364 5468 3672 5477
rect 3364 5466 3370 5468
rect 3426 5466 3450 5468
rect 3506 5466 3530 5468
rect 3586 5466 3610 5468
rect 3666 5466 3672 5468
rect 3426 5414 3428 5466
rect 3608 5414 3610 5466
rect 3364 5412 3370 5414
rect 3426 5412 3450 5414
rect 3506 5412 3530 5414
rect 3586 5412 3610 5414
rect 3666 5412 3672 5414
rect 3364 5403 3672 5412
rect 3988 5370 4016 5646
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3252 3534 3280 5102
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 4826 3740 4966
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3364 4380 3672 4389
rect 3364 4378 3370 4380
rect 3426 4378 3450 4380
rect 3506 4378 3530 4380
rect 3586 4378 3610 4380
rect 3666 4378 3672 4380
rect 3426 4326 3428 4378
rect 3608 4326 3610 4378
rect 3364 4324 3370 4326
rect 3426 4324 3450 4326
rect 3506 4324 3530 4326
rect 3586 4324 3610 4326
rect 3666 4324 3672 4326
rect 3364 4315 3672 4324
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3738 3372 4082
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3252 2922 3280 3470
rect 3364 3292 3672 3301
rect 3364 3290 3370 3292
rect 3426 3290 3450 3292
rect 3506 3290 3530 3292
rect 3586 3290 3610 3292
rect 3666 3290 3672 3292
rect 3426 3238 3428 3290
rect 3608 3238 3610 3290
rect 3364 3236 3370 3238
rect 3426 3236 3450 3238
rect 3506 3236 3530 3238
rect 3586 3236 3610 3238
rect 3666 3236 3672 3238
rect 3364 3227 3672 3236
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3712 2854 3740 3470
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 2157 2748 2465 2757
rect 2157 2746 2163 2748
rect 2219 2746 2243 2748
rect 2299 2746 2323 2748
rect 2379 2746 2403 2748
rect 2459 2746 2465 2748
rect 2219 2694 2221 2746
rect 2401 2694 2403 2746
rect 2157 2692 2163 2694
rect 2219 2692 2243 2694
rect 2299 2692 2323 2694
rect 2379 2692 2403 2694
rect 2459 2692 2465 2694
rect 2157 2683 2465 2692
rect 2884 2746 3188 2774
rect 2884 2650 2912 2746
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3712 2514 3740 2790
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2976 800 3004 2382
rect 3988 2378 4016 4014
rect 4066 3496 4122 3505
rect 4172 3482 4200 6666
rect 5644 6322 5672 7346
rect 6196 6662 6224 7754
rect 6380 7750 6408 8366
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8022 6868 8230
rect 6987 8188 7295 8197
rect 6987 8186 6993 8188
rect 7049 8186 7073 8188
rect 7129 8186 7153 8188
rect 7209 8186 7233 8188
rect 7289 8186 7295 8188
rect 7049 8134 7051 8186
rect 7231 8134 7233 8186
rect 6987 8132 6993 8134
rect 7049 8132 7073 8134
rect 7129 8132 7153 8134
rect 7209 8132 7233 8134
rect 7289 8132 7295 8134
rect 6987 8123 7295 8132
rect 7484 8090 7512 9522
rect 7576 8906 7604 9658
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7668 8634 7696 9930
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9586 7788 9862
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7852 9110 7880 10542
rect 7944 10198 7972 10950
rect 8194 10908 8502 10917
rect 8194 10906 8200 10908
rect 8256 10906 8280 10908
rect 8336 10906 8360 10908
rect 8416 10906 8440 10908
rect 8496 10906 8502 10908
rect 8256 10854 8258 10906
rect 8438 10854 8440 10906
rect 8194 10852 8200 10854
rect 8256 10852 8280 10854
rect 8336 10852 8360 10854
rect 8416 10852 8440 10854
rect 8496 10852 8502 10854
rect 8194 10843 8502 10852
rect 9140 10810 9168 11018
rect 10609 10908 10917 10917
rect 10609 10906 10615 10908
rect 10671 10906 10695 10908
rect 10751 10906 10775 10908
rect 10831 10906 10855 10908
rect 10911 10906 10917 10908
rect 10671 10854 10673 10906
rect 10853 10854 10855 10906
rect 10609 10852 10615 10854
rect 10671 10852 10695 10854
rect 10751 10852 10775 10854
rect 10831 10852 10855 10854
rect 10911 10852 10917 10854
rect 10609 10843 10917 10852
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8128 10198 8156 10746
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8404 10266 8432 10678
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7944 9382 7972 10134
rect 8128 9722 8156 10134
rect 8220 10062 8248 10202
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8194 9820 8502 9829
rect 8194 9818 8200 9820
rect 8256 9818 8280 9820
rect 8336 9818 8360 9820
rect 8416 9818 8440 9820
rect 8496 9818 8502 9820
rect 8256 9766 8258 9818
rect 8438 9766 8440 9818
rect 8194 9764 8200 9766
rect 8256 9764 8280 9766
rect 8336 9764 8360 9766
rect 8416 9764 8440 9766
rect 8496 9764 8502 9766
rect 8194 9755 8502 9764
rect 8680 9722 8708 10066
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7944 8906 7972 9318
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7410 6408 7686
rect 7484 7546 7512 8026
rect 7760 7970 7788 8842
rect 7944 8514 7972 8842
rect 8036 8634 8064 8842
rect 8128 8634 8156 9318
rect 8194 8732 8502 8741
rect 8194 8730 8200 8732
rect 8256 8730 8280 8732
rect 8336 8730 8360 8732
rect 8416 8730 8440 8732
rect 8496 8730 8502 8732
rect 8256 8678 8258 8730
rect 8438 8678 8440 8730
rect 8194 8676 8200 8678
rect 8256 8676 8280 8678
rect 8336 8676 8360 8678
rect 8416 8676 8440 8678
rect 8496 8676 8502 8678
rect 8194 8667 8502 8676
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7944 8486 8064 8514
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7576 7942 7788 7970
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6987 7100 7295 7109
rect 6987 7098 6993 7100
rect 7049 7098 7073 7100
rect 7129 7098 7153 7100
rect 7209 7098 7233 7100
rect 7289 7098 7295 7100
rect 7049 7046 7051 7098
rect 7231 7046 7233 7098
rect 6987 7044 6993 7046
rect 7049 7044 7073 7046
rect 7129 7044 7153 7046
rect 7209 7044 7233 7046
rect 7289 7044 7295 7046
rect 6987 7035 7295 7044
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5779 6556 6087 6565
rect 5779 6554 5785 6556
rect 5841 6554 5865 6556
rect 5921 6554 5945 6556
rect 6001 6554 6025 6556
rect 6081 6554 6087 6556
rect 5841 6502 5843 6554
rect 6023 6502 6025 6554
rect 5779 6500 5785 6502
rect 5841 6500 5865 6502
rect 5921 6500 5945 6502
rect 6001 6500 6025 6502
rect 6081 6500 6087 6502
rect 5779 6491 6087 6500
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 4572 6012 4880 6021
rect 4572 6010 4578 6012
rect 4634 6010 4658 6012
rect 4714 6010 4738 6012
rect 4794 6010 4818 6012
rect 4874 6010 4880 6012
rect 4634 5958 4636 6010
rect 4816 5958 4818 6010
rect 4572 5956 4578 5958
rect 4634 5956 4658 5958
rect 4714 5956 4738 5958
rect 4794 5956 4818 5958
rect 4874 5956 4880 5958
rect 4572 5947 4880 5956
rect 5276 5574 5304 6258
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4724 5370 4752 5510
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4572 4924 4880 4933
rect 4572 4922 4578 4924
rect 4634 4922 4658 4924
rect 4714 4922 4738 4924
rect 4794 4922 4818 4924
rect 4874 4922 4880 4924
rect 4634 4870 4636 4922
rect 4816 4870 4818 4922
rect 4572 4868 4578 4870
rect 4634 4868 4658 4870
rect 4714 4868 4738 4870
rect 4794 4868 4818 4870
rect 4874 4868 4880 4870
rect 4572 4859 4880 4868
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4078 4476 4422
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 5276 4010 5304 5510
rect 5552 5302 5580 6054
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5644 5030 5672 5510
rect 5779 5468 6087 5477
rect 5779 5466 5785 5468
rect 5841 5466 5865 5468
rect 5921 5466 5945 5468
rect 6001 5466 6025 5468
rect 6081 5466 6087 5468
rect 5841 5414 5843 5466
rect 6023 5414 6025 5466
rect 5779 5412 5785 5414
rect 5841 5412 5865 5414
rect 5921 5412 5945 5414
rect 6001 5412 6025 5414
rect 6081 5412 6087 5414
rect 5779 5403 6087 5412
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 4572 3836 4880 3845
rect 4572 3834 4578 3836
rect 4634 3834 4658 3836
rect 4714 3834 4738 3836
rect 4794 3834 4818 3836
rect 4874 3834 4880 3836
rect 4634 3782 4636 3834
rect 4816 3782 4818 3834
rect 4572 3780 4578 3782
rect 4634 3780 4658 3782
rect 4714 3780 4738 3782
rect 4794 3780 4818 3782
rect 4874 3780 4880 3782
rect 4572 3771 4880 3780
rect 4122 3454 4200 3482
rect 5448 3460 5500 3466
rect 4066 3431 4122 3440
rect 5448 3402 5500 3408
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 2774 4108 2858
rect 4080 2746 4200 2774
rect 4172 2378 4200 2746
rect 4572 2748 4880 2757
rect 4572 2746 4578 2748
rect 4634 2746 4658 2748
rect 4714 2746 4738 2748
rect 4794 2746 4818 2748
rect 4874 2746 4880 2748
rect 4634 2694 4636 2746
rect 4816 2694 4818 2746
rect 4572 2692 4578 2694
rect 4634 2692 4658 2694
rect 4714 2692 4738 2694
rect 4794 2692 4818 2694
rect 4874 2692 4880 2694
rect 4572 2683 4880 2692
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 5460 2310 5488 3402
rect 5552 3398 5580 4082
rect 5644 3602 5672 4966
rect 5779 4380 6087 4389
rect 5779 4378 5785 4380
rect 5841 4378 5865 4380
rect 5921 4378 5945 4380
rect 6001 4378 6025 4380
rect 6081 4378 6087 4380
rect 5841 4326 5843 4378
rect 6023 4326 6025 4378
rect 5779 4324 5785 4326
rect 5841 4324 5865 4326
rect 5921 4324 5945 4326
rect 6001 4324 6025 4326
rect 6081 4324 6087 4326
rect 5779 4315 6087 4324
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3738 5764 3878
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 2990 5580 3334
rect 5779 3292 6087 3301
rect 5779 3290 5785 3292
rect 5841 3290 5865 3292
rect 5921 3290 5945 3292
rect 6001 3290 6025 3292
rect 6081 3290 6087 3292
rect 5841 3238 5843 3290
rect 6023 3238 6025 3290
rect 5779 3236 5785 3238
rect 5841 3236 5865 3238
rect 5921 3236 5945 3238
rect 6001 3236 6025 3238
rect 6081 3236 6087 3238
rect 5779 3227 6087 3236
rect 6196 3126 6224 6598
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5642 6316 6054
rect 6987 6012 7295 6021
rect 6987 6010 6993 6012
rect 7049 6010 7073 6012
rect 7129 6010 7153 6012
rect 7209 6010 7233 6012
rect 7289 6010 7295 6012
rect 7049 5958 7051 6010
rect 7231 5958 7233 6010
rect 6987 5956 6993 5958
rect 7049 5956 7073 5958
rect 7129 5956 7153 5958
rect 7209 5956 7233 5958
rect 7289 5956 7295 5958
rect 6987 5947 7295 5956
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6288 5370 6316 5578
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6288 3398 6316 5306
rect 6987 4924 7295 4933
rect 6987 4922 6993 4924
rect 7049 4922 7073 4924
rect 7129 4922 7153 4924
rect 7209 4922 7233 4924
rect 7289 4922 7295 4924
rect 7049 4870 7051 4922
rect 7231 4870 7233 4922
rect 6987 4868 6993 4870
rect 7049 4868 7073 4870
rect 7129 4868 7153 4870
rect 7209 4868 7233 4870
rect 7289 4868 7295 4870
rect 6987 4859 7295 4868
rect 7576 4758 7604 7942
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7546 7788 7822
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7852 7342 7880 8298
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7760 6458 7788 6666
rect 7944 6458 7972 7686
rect 8036 7478 8064 8486
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8194 7644 8502 7653
rect 8194 7642 8200 7644
rect 8256 7642 8280 7644
rect 8336 7642 8360 7644
rect 8416 7642 8440 7644
rect 8496 7642 8502 7644
rect 8256 7590 8258 7642
rect 8438 7590 8440 7642
rect 8194 7588 8200 7590
rect 8256 7588 8280 7590
rect 8336 7588 8360 7590
rect 8416 7588 8440 7590
rect 8496 7588 8502 7590
rect 8194 7579 8502 7588
rect 8588 7546 8616 7822
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 7002 8616 7278
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8194 6556 8502 6565
rect 8194 6554 8200 6556
rect 8256 6554 8280 6556
rect 8336 6554 8360 6556
rect 8416 6554 8440 6556
rect 8496 6554 8502 6556
rect 8256 6502 8258 6554
rect 8438 6502 8440 6554
rect 8194 6500 8200 6502
rect 8256 6500 8280 6502
rect 8336 6500 8360 6502
rect 8416 6500 8440 6502
rect 8496 6500 8502 6502
rect 8194 6491 8502 6500
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8588 6118 8616 6598
rect 8680 6322 8708 7210
rect 8864 6746 8892 10610
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 9220 10464 9272 10470
rect 10888 10441 10916 10474
rect 9220 10406 9272 10412
rect 10874 10432 10930 10441
rect 9232 10130 9260 10406
rect 9402 10364 9710 10373
rect 10874 10367 10930 10376
rect 9402 10362 9408 10364
rect 9464 10362 9488 10364
rect 9544 10362 9568 10364
rect 9624 10362 9648 10364
rect 9704 10362 9710 10364
rect 9464 10310 9466 10362
rect 9646 10310 9648 10362
rect 9402 10308 9408 10310
rect 9464 10308 9488 10310
rect 9544 10308 9568 10310
rect 9624 10308 9648 10310
rect 9704 10308 9710 10310
rect 9402 10299 9710 10308
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9654 9536 9862
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9402 9276 9710 9285
rect 9402 9274 9408 9276
rect 9464 9274 9488 9276
rect 9544 9274 9568 9276
rect 9624 9274 9648 9276
rect 9704 9274 9710 9276
rect 9464 9222 9466 9274
rect 9646 9222 9648 9274
rect 9402 9220 9408 9222
rect 9464 9220 9488 9222
rect 9544 9220 9568 9222
rect 9624 9220 9648 9222
rect 9704 9220 9710 9222
rect 9402 9211 9710 9220
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7546 8984 7686
rect 9140 7546 9168 7958
rect 9232 7546 9260 8774
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7886 9352 8230
rect 9402 8188 9710 8197
rect 9402 8186 9408 8188
rect 9464 8186 9488 8188
rect 9544 8186 9568 8188
rect 9624 8186 9648 8188
rect 9704 8186 9710 8188
rect 9464 8134 9466 8186
rect 9646 8134 9648 8186
rect 9402 8132 9408 8134
rect 9464 8132 9488 8134
rect 9544 8132 9568 8134
rect 9624 8132 9648 8134
rect 9704 8132 9710 8134
rect 9402 8123 9710 8132
rect 9876 8090 9904 8842
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9956 7880 10008 7886
rect 10008 7828 10088 7834
rect 9956 7822 10088 7828
rect 9968 7806 10088 7822
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 6934 9352 7346
rect 9402 7100 9710 7109
rect 9402 7098 9408 7100
rect 9464 7098 9488 7100
rect 9544 7098 9568 7100
rect 9624 7098 9648 7100
rect 9704 7098 9710 7100
rect 9464 7046 9466 7098
rect 9646 7046 9648 7098
rect 9402 7044 9408 7046
rect 9464 7044 9488 7046
rect 9544 7044 9568 7046
rect 9624 7044 9648 7046
rect 9704 7044 9710 7046
rect 9402 7035 9710 7044
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 8864 6718 8984 6746
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6458 8892 6598
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7576 4146 7604 4694
rect 7668 4146 7696 5850
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 6987 3836 7295 3845
rect 6987 3834 6993 3836
rect 7049 3834 7073 3836
rect 7129 3834 7153 3836
rect 7209 3834 7233 3836
rect 7289 3834 7295 3836
rect 7049 3782 7051 3834
rect 7231 3782 7233 3834
rect 6987 3780 6993 3782
rect 7049 3780 7073 3782
rect 7129 3780 7153 3782
rect 7209 3780 7233 3782
rect 7289 3780 7295 3782
rect 6987 3771 7295 3780
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7300 3126 7328 3334
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5552 2650 5580 2926
rect 7576 2922 7604 4082
rect 7760 3738 7788 4082
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7852 3194 7880 5510
rect 8194 5468 8502 5477
rect 8194 5466 8200 5468
rect 8256 5466 8280 5468
rect 8336 5466 8360 5468
rect 8416 5466 8440 5468
rect 8496 5466 8502 5468
rect 8256 5414 8258 5466
rect 8438 5414 8440 5466
rect 8194 5412 8200 5414
rect 8256 5412 8280 5414
rect 8336 5412 8360 5414
rect 8416 5412 8440 5414
rect 8496 5412 8502 5414
rect 8194 5403 8502 5412
rect 8588 5234 8616 6054
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7944 3466 7972 4422
rect 8036 4146 8064 4422
rect 8194 4380 8502 4389
rect 8194 4378 8200 4380
rect 8256 4378 8280 4380
rect 8336 4378 8360 4380
rect 8416 4378 8440 4380
rect 8496 4378 8502 4380
rect 8256 4326 8258 4378
rect 8438 4326 8440 4378
rect 8194 4324 8200 4326
rect 8256 4324 8280 4326
rect 8336 4324 8360 4326
rect 8416 4324 8440 4326
rect 8496 4324 8502 4326
rect 8194 4315 8502 4324
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8220 3534 8248 3946
rect 8588 3602 8616 5170
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4026 8708 4626
rect 8772 4146 8800 4966
rect 8864 4758 8892 5850
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8852 4072 8904 4078
rect 8680 4020 8852 4026
rect 8680 4014 8904 4020
rect 8680 3998 8892 4014
rect 8680 3738 8708 3998
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8208 3528 8260 3534
rect 8128 3476 8208 3482
rect 8128 3470 8260 3476
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 8128 3454 8248 3470
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 6987 2748 7295 2757
rect 6987 2746 6993 2748
rect 7049 2746 7073 2748
rect 7129 2746 7153 2748
rect 7209 2746 7233 2748
rect 7289 2746 7295 2748
rect 7049 2694 7051 2746
rect 7231 2694 7233 2746
rect 6987 2692 6993 2694
rect 7049 2692 7073 2694
rect 7129 2692 7153 2694
rect 7209 2692 7233 2694
rect 7289 2692 7295 2694
rect 6987 2683 7295 2692
rect 7576 2650 7604 2858
rect 7944 2650 7972 2994
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8128 2446 8156 3454
rect 8194 3292 8502 3301
rect 8194 3290 8200 3292
rect 8256 3290 8280 3292
rect 8336 3290 8360 3292
rect 8416 3290 8440 3292
rect 8496 3290 8502 3292
rect 8256 3238 8258 3290
rect 8438 3238 8440 3290
rect 8194 3236 8200 3238
rect 8256 3236 8280 3238
rect 8336 3236 8360 3238
rect 8416 3236 8440 3238
rect 8496 3236 8502 3238
rect 8194 3227 8502 3236
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 2582 8432 3130
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 3364 2204 3672 2213
rect 3364 2202 3370 2204
rect 3426 2202 3450 2204
rect 3506 2202 3530 2204
rect 3586 2202 3610 2204
rect 3666 2202 3672 2204
rect 3426 2150 3428 2202
rect 3608 2150 3610 2202
rect 3364 2148 3370 2150
rect 3426 2148 3450 2150
rect 3506 2148 3530 2150
rect 3586 2148 3610 2150
rect 3666 2148 3672 2150
rect 3364 2139 3672 2148
rect 5779 2204 6087 2213
rect 5779 2202 5785 2204
rect 5841 2202 5865 2204
rect 5921 2202 5945 2204
rect 6001 2202 6025 2204
rect 6081 2202 6087 2204
rect 5841 2150 5843 2202
rect 6023 2150 6025 2202
rect 5779 2148 5785 2150
rect 5841 2148 5865 2150
rect 5921 2148 5945 2150
rect 6001 2148 6025 2150
rect 6081 2148 6087 2150
rect 5779 2139 6087 2148
rect 8194 2204 8502 2213
rect 8194 2202 8200 2204
rect 8256 2202 8280 2204
rect 8336 2202 8360 2204
rect 8416 2202 8440 2204
rect 8496 2202 8502 2204
rect 8256 2150 8258 2202
rect 8438 2150 8440 2202
rect 8194 2148 8200 2150
rect 8256 2148 8280 2150
rect 8336 2148 8360 2150
rect 8416 2148 8440 2150
rect 8496 2148 8502 2150
rect 8194 2139 8502 2148
rect 8772 1306 8800 2314
rect 8956 2310 8984 6718
rect 9402 6012 9710 6021
rect 9402 6010 9408 6012
rect 9464 6010 9488 6012
rect 9544 6010 9568 6012
rect 9624 6010 9648 6012
rect 9704 6010 9710 6012
rect 9464 5958 9466 6010
rect 9646 5958 9648 6010
rect 9402 5956 9408 5958
rect 9464 5956 9488 5958
rect 9544 5956 9568 5958
rect 9624 5956 9648 5958
rect 9704 5956 9710 5958
rect 9402 5947 9710 5956
rect 9784 5914 9812 7686
rect 9968 7206 9996 7686
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9876 6866 9904 7142
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9968 5710 9996 7142
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9048 4622 9076 5510
rect 9232 5302 9260 5510
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4690 9168 4966
rect 9402 4924 9710 4933
rect 9402 4922 9408 4924
rect 9464 4922 9488 4924
rect 9544 4922 9568 4924
rect 9624 4922 9648 4924
rect 9704 4922 9710 4924
rect 9464 4870 9466 4922
rect 9646 4870 9648 4922
rect 9402 4868 9408 4870
rect 9464 4868 9488 4870
rect 9544 4868 9568 4870
rect 9624 4868 9648 4870
rect 9704 4868 9710 4870
rect 9402 4859 9710 4868
rect 9784 4826 9812 5646
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4690 9904 4966
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9048 3194 9076 4014
rect 9140 3534 9168 4626
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 3942 9260 4558
rect 9876 4146 9904 4626
rect 10060 4146 10088 7806
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10152 5710 10180 7686
rect 10244 7410 10272 7686
rect 10336 7478 10364 7686
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 6458 10272 7346
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9402 3836 9710 3845
rect 9402 3834 9408 3836
rect 9464 3834 9488 3836
rect 9544 3834 9568 3836
rect 9624 3834 9648 3836
rect 9704 3834 9710 3836
rect 9464 3782 9466 3834
rect 9646 3782 9648 3834
rect 9402 3780 9408 3782
rect 9464 3780 9488 3782
rect 9544 3780 9568 3782
rect 9624 3780 9648 3782
rect 9704 3780 9710 3782
rect 9402 3771 9710 3780
rect 9968 3738 9996 4014
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 3194 9904 3402
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9048 2514 9076 3130
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9402 2748 9710 2757
rect 9402 2746 9408 2748
rect 9464 2746 9488 2748
rect 9544 2746 9568 2748
rect 9624 2746 9648 2748
rect 9704 2746 9710 2748
rect 9464 2694 9466 2746
rect 9646 2694 9648 2746
rect 9402 2692 9408 2694
rect 9464 2692 9488 2694
rect 9544 2692 9568 2694
rect 9624 2692 9648 2694
rect 9704 2692 9710 2694
rect 9402 2683 9710 2692
rect 9784 2650 9812 2790
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10336 2514 10364 3674
rect 10428 3194 10456 10202
rect 10609 9820 10917 9829
rect 10609 9818 10615 9820
rect 10671 9818 10695 9820
rect 10751 9818 10775 9820
rect 10831 9818 10855 9820
rect 10911 9818 10917 9820
rect 10671 9766 10673 9818
rect 10853 9766 10855 9818
rect 10609 9764 10615 9766
rect 10671 9764 10695 9766
rect 10751 9764 10775 9766
rect 10831 9764 10855 9766
rect 10911 9764 10917 9766
rect 10609 9755 10917 9764
rect 10609 8732 10917 8741
rect 10609 8730 10615 8732
rect 10671 8730 10695 8732
rect 10751 8730 10775 8732
rect 10831 8730 10855 8732
rect 10911 8730 10917 8732
rect 10671 8678 10673 8730
rect 10853 8678 10855 8730
rect 10609 8676 10615 8678
rect 10671 8676 10695 8678
rect 10751 8676 10775 8678
rect 10831 8676 10855 8678
rect 10911 8676 10917 8678
rect 10609 8667 10917 8676
rect 10609 7644 10917 7653
rect 10609 7642 10615 7644
rect 10671 7642 10695 7644
rect 10751 7642 10775 7644
rect 10831 7642 10855 7644
rect 10911 7642 10917 7644
rect 10671 7590 10673 7642
rect 10853 7590 10855 7642
rect 10609 7588 10615 7590
rect 10671 7588 10695 7590
rect 10751 7588 10775 7590
rect 10831 7588 10855 7590
rect 10911 7588 10917 7590
rect 10609 7579 10917 7588
rect 10609 6556 10917 6565
rect 10609 6554 10615 6556
rect 10671 6554 10695 6556
rect 10751 6554 10775 6556
rect 10831 6554 10855 6556
rect 10911 6554 10917 6556
rect 10671 6502 10673 6554
rect 10853 6502 10855 6554
rect 10609 6500 10615 6502
rect 10671 6500 10695 6502
rect 10751 6500 10775 6502
rect 10831 6500 10855 6502
rect 10911 6500 10917 6502
rect 10609 6491 10917 6500
rect 10609 5468 10917 5477
rect 10609 5466 10615 5468
rect 10671 5466 10695 5468
rect 10751 5466 10775 5468
rect 10831 5466 10855 5468
rect 10911 5466 10917 5468
rect 10671 5414 10673 5466
rect 10853 5414 10855 5466
rect 10609 5412 10615 5414
rect 10671 5412 10695 5414
rect 10751 5412 10775 5414
rect 10831 5412 10855 5414
rect 10911 5412 10917 5414
rect 10609 5403 10917 5412
rect 10609 4380 10917 4389
rect 10609 4378 10615 4380
rect 10671 4378 10695 4380
rect 10751 4378 10775 4380
rect 10831 4378 10855 4380
rect 10911 4378 10917 4380
rect 10671 4326 10673 4378
rect 10853 4326 10855 4378
rect 10609 4324 10615 4326
rect 10671 4324 10695 4326
rect 10751 4324 10775 4326
rect 10831 4324 10855 4326
rect 10911 4324 10917 4326
rect 10609 4315 10917 4324
rect 10609 3292 10917 3301
rect 10609 3290 10615 3292
rect 10671 3290 10695 3292
rect 10751 3290 10775 3292
rect 10831 3290 10855 3292
rect 10911 3290 10917 3292
rect 10671 3238 10673 3290
rect 10853 3238 10855 3290
rect 10609 3236 10615 3238
rect 10671 3236 10695 3238
rect 10751 3236 10775 3238
rect 10831 3236 10855 3238
rect 10911 3236 10917 3238
rect 10609 3227 10917 3236
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10874 3088 10930 3097
rect 10874 3023 10876 3032
rect 10928 3023 10930 3032
rect 10876 2994 10928 3000
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 10609 2204 10917 2213
rect 10609 2202 10615 2204
rect 10671 2202 10695 2204
rect 10751 2202 10775 2204
rect 10831 2202 10855 2204
rect 10911 2202 10917 2204
rect 10671 2150 10673 2202
rect 10853 2150 10855 2202
rect 10609 2148 10615 2150
rect 10671 2148 10695 2150
rect 10751 2148 10775 2150
rect 10831 2148 10855 2150
rect 10911 2148 10917 2150
rect 10609 2139 10917 2148
rect 8772 1278 8984 1306
rect 8956 800 8984 1278
rect 2962 0 3018 800
rect 8942 0 8998 800
<< via2 >>
rect 2163 11450 2219 11452
rect 2243 11450 2299 11452
rect 2323 11450 2379 11452
rect 2403 11450 2459 11452
rect 2163 11398 2209 11450
rect 2209 11398 2219 11450
rect 2243 11398 2273 11450
rect 2273 11398 2285 11450
rect 2285 11398 2299 11450
rect 2323 11398 2337 11450
rect 2337 11398 2349 11450
rect 2349 11398 2379 11450
rect 2403 11398 2413 11450
rect 2413 11398 2459 11450
rect 2163 11396 2219 11398
rect 2243 11396 2299 11398
rect 2323 11396 2379 11398
rect 2403 11396 2459 11398
rect 4578 11450 4634 11452
rect 4658 11450 4714 11452
rect 4738 11450 4794 11452
rect 4818 11450 4874 11452
rect 4578 11398 4624 11450
rect 4624 11398 4634 11450
rect 4658 11398 4688 11450
rect 4688 11398 4700 11450
rect 4700 11398 4714 11450
rect 4738 11398 4752 11450
rect 4752 11398 4764 11450
rect 4764 11398 4794 11450
rect 4818 11398 4828 11450
rect 4828 11398 4874 11450
rect 4578 11396 4634 11398
rect 4658 11396 4714 11398
rect 4738 11396 4794 11398
rect 4818 11396 4874 11398
rect 6993 11450 7049 11452
rect 7073 11450 7129 11452
rect 7153 11450 7209 11452
rect 7233 11450 7289 11452
rect 6993 11398 7039 11450
rect 7039 11398 7049 11450
rect 7073 11398 7103 11450
rect 7103 11398 7115 11450
rect 7115 11398 7129 11450
rect 7153 11398 7167 11450
rect 7167 11398 7179 11450
rect 7179 11398 7209 11450
rect 7233 11398 7243 11450
rect 7243 11398 7289 11450
rect 6993 11396 7049 11398
rect 7073 11396 7129 11398
rect 7153 11396 7209 11398
rect 7233 11396 7289 11398
rect 9408 11450 9464 11452
rect 9488 11450 9544 11452
rect 9568 11450 9624 11452
rect 9648 11450 9704 11452
rect 9408 11398 9454 11450
rect 9454 11398 9464 11450
rect 9488 11398 9518 11450
rect 9518 11398 9530 11450
rect 9530 11398 9544 11450
rect 9568 11398 9582 11450
rect 9582 11398 9594 11450
rect 9594 11398 9624 11450
rect 9648 11398 9658 11450
rect 9658 11398 9704 11450
rect 9408 11396 9464 11398
rect 9488 11396 9544 11398
rect 9568 11396 9624 11398
rect 9648 11396 9704 11398
rect 938 10376 994 10432
rect 2163 10362 2219 10364
rect 2243 10362 2299 10364
rect 2323 10362 2379 10364
rect 2403 10362 2459 10364
rect 2163 10310 2209 10362
rect 2209 10310 2219 10362
rect 2243 10310 2273 10362
rect 2273 10310 2285 10362
rect 2285 10310 2299 10362
rect 2323 10310 2337 10362
rect 2337 10310 2349 10362
rect 2349 10310 2379 10362
rect 2403 10310 2413 10362
rect 2413 10310 2459 10362
rect 2163 10308 2219 10310
rect 2243 10308 2299 10310
rect 2323 10308 2379 10310
rect 2403 10308 2459 10310
rect 2163 9274 2219 9276
rect 2243 9274 2299 9276
rect 2323 9274 2379 9276
rect 2403 9274 2459 9276
rect 2163 9222 2209 9274
rect 2209 9222 2219 9274
rect 2243 9222 2273 9274
rect 2273 9222 2285 9274
rect 2285 9222 2299 9274
rect 2323 9222 2337 9274
rect 2337 9222 2349 9274
rect 2349 9222 2379 9274
rect 2403 9222 2413 9274
rect 2413 9222 2459 9274
rect 2163 9220 2219 9222
rect 2243 9220 2299 9222
rect 2323 9220 2379 9222
rect 2403 9220 2459 9222
rect 2163 8186 2219 8188
rect 2243 8186 2299 8188
rect 2323 8186 2379 8188
rect 2403 8186 2459 8188
rect 2163 8134 2209 8186
rect 2209 8134 2219 8186
rect 2243 8134 2273 8186
rect 2273 8134 2285 8186
rect 2285 8134 2299 8186
rect 2323 8134 2337 8186
rect 2337 8134 2349 8186
rect 2349 8134 2379 8186
rect 2403 8134 2413 8186
rect 2413 8134 2459 8186
rect 2163 8132 2219 8134
rect 2243 8132 2299 8134
rect 2323 8132 2379 8134
rect 2403 8132 2459 8134
rect 2163 7098 2219 7100
rect 2243 7098 2299 7100
rect 2323 7098 2379 7100
rect 2403 7098 2459 7100
rect 2163 7046 2209 7098
rect 2209 7046 2219 7098
rect 2243 7046 2273 7098
rect 2273 7046 2285 7098
rect 2285 7046 2299 7098
rect 2323 7046 2337 7098
rect 2337 7046 2349 7098
rect 2349 7046 2379 7098
rect 2403 7046 2413 7098
rect 2413 7046 2459 7098
rect 2163 7044 2219 7046
rect 2243 7044 2299 7046
rect 2323 7044 2379 7046
rect 2403 7044 2459 7046
rect 3370 10906 3426 10908
rect 3450 10906 3506 10908
rect 3530 10906 3586 10908
rect 3610 10906 3666 10908
rect 3370 10854 3416 10906
rect 3416 10854 3426 10906
rect 3450 10854 3480 10906
rect 3480 10854 3492 10906
rect 3492 10854 3506 10906
rect 3530 10854 3544 10906
rect 3544 10854 3556 10906
rect 3556 10854 3586 10906
rect 3610 10854 3620 10906
rect 3620 10854 3666 10906
rect 3370 10852 3426 10854
rect 3450 10852 3506 10854
rect 3530 10852 3586 10854
rect 3610 10852 3666 10854
rect 5785 10906 5841 10908
rect 5865 10906 5921 10908
rect 5945 10906 6001 10908
rect 6025 10906 6081 10908
rect 5785 10854 5831 10906
rect 5831 10854 5841 10906
rect 5865 10854 5895 10906
rect 5895 10854 5907 10906
rect 5907 10854 5921 10906
rect 5945 10854 5959 10906
rect 5959 10854 5971 10906
rect 5971 10854 6001 10906
rect 6025 10854 6035 10906
rect 6035 10854 6081 10906
rect 5785 10852 5841 10854
rect 5865 10852 5921 10854
rect 5945 10852 6001 10854
rect 6025 10852 6081 10854
rect 3370 9818 3426 9820
rect 3450 9818 3506 9820
rect 3530 9818 3586 9820
rect 3610 9818 3666 9820
rect 3370 9766 3416 9818
rect 3416 9766 3426 9818
rect 3450 9766 3480 9818
rect 3480 9766 3492 9818
rect 3492 9766 3506 9818
rect 3530 9766 3544 9818
rect 3544 9766 3556 9818
rect 3556 9766 3586 9818
rect 3610 9766 3620 9818
rect 3620 9766 3666 9818
rect 3370 9764 3426 9766
rect 3450 9764 3506 9766
rect 3530 9764 3586 9766
rect 3610 9764 3666 9766
rect 3370 8730 3426 8732
rect 3450 8730 3506 8732
rect 3530 8730 3586 8732
rect 3610 8730 3666 8732
rect 3370 8678 3416 8730
rect 3416 8678 3426 8730
rect 3450 8678 3480 8730
rect 3480 8678 3492 8730
rect 3492 8678 3506 8730
rect 3530 8678 3544 8730
rect 3544 8678 3556 8730
rect 3556 8678 3586 8730
rect 3610 8678 3620 8730
rect 3620 8678 3666 8730
rect 3370 8676 3426 8678
rect 3450 8676 3506 8678
rect 3530 8676 3586 8678
rect 3610 8676 3666 8678
rect 2163 6010 2219 6012
rect 2243 6010 2299 6012
rect 2323 6010 2379 6012
rect 2403 6010 2459 6012
rect 2163 5958 2209 6010
rect 2209 5958 2219 6010
rect 2243 5958 2273 6010
rect 2273 5958 2285 6010
rect 2285 5958 2299 6010
rect 2323 5958 2337 6010
rect 2337 5958 2349 6010
rect 2349 5958 2379 6010
rect 2403 5958 2413 6010
rect 2413 5958 2459 6010
rect 2163 5956 2219 5958
rect 2243 5956 2299 5958
rect 2323 5956 2379 5958
rect 2403 5956 2459 5958
rect 2163 4922 2219 4924
rect 2243 4922 2299 4924
rect 2323 4922 2379 4924
rect 2403 4922 2459 4924
rect 2163 4870 2209 4922
rect 2209 4870 2219 4922
rect 2243 4870 2273 4922
rect 2273 4870 2285 4922
rect 2285 4870 2299 4922
rect 2323 4870 2337 4922
rect 2337 4870 2349 4922
rect 2349 4870 2379 4922
rect 2403 4870 2413 4922
rect 2413 4870 2459 4922
rect 2163 4868 2219 4870
rect 2243 4868 2299 4870
rect 2323 4868 2379 4870
rect 2403 4868 2459 4870
rect 2163 3834 2219 3836
rect 2243 3834 2299 3836
rect 2323 3834 2379 3836
rect 2403 3834 2459 3836
rect 2163 3782 2209 3834
rect 2209 3782 2219 3834
rect 2243 3782 2273 3834
rect 2273 3782 2285 3834
rect 2285 3782 2299 3834
rect 2323 3782 2337 3834
rect 2337 3782 2349 3834
rect 2349 3782 2379 3834
rect 2403 3782 2413 3834
rect 2413 3782 2459 3834
rect 2163 3780 2219 3782
rect 2243 3780 2299 3782
rect 2323 3780 2379 3782
rect 2403 3780 2459 3782
rect 3370 7642 3426 7644
rect 3450 7642 3506 7644
rect 3530 7642 3586 7644
rect 3610 7642 3666 7644
rect 3370 7590 3416 7642
rect 3416 7590 3426 7642
rect 3450 7590 3480 7642
rect 3480 7590 3492 7642
rect 3492 7590 3506 7642
rect 3530 7590 3544 7642
rect 3544 7590 3556 7642
rect 3556 7590 3586 7642
rect 3610 7590 3620 7642
rect 3620 7590 3666 7642
rect 3370 7588 3426 7590
rect 3450 7588 3506 7590
rect 3530 7588 3586 7590
rect 3610 7588 3666 7590
rect 4578 10362 4634 10364
rect 4658 10362 4714 10364
rect 4738 10362 4794 10364
rect 4818 10362 4874 10364
rect 4578 10310 4624 10362
rect 4624 10310 4634 10362
rect 4658 10310 4688 10362
rect 4688 10310 4700 10362
rect 4700 10310 4714 10362
rect 4738 10310 4752 10362
rect 4752 10310 4764 10362
rect 4764 10310 4794 10362
rect 4818 10310 4828 10362
rect 4828 10310 4874 10362
rect 4578 10308 4634 10310
rect 4658 10308 4714 10310
rect 4738 10308 4794 10310
rect 4818 10308 4874 10310
rect 4578 9274 4634 9276
rect 4658 9274 4714 9276
rect 4738 9274 4794 9276
rect 4818 9274 4874 9276
rect 4578 9222 4624 9274
rect 4624 9222 4634 9274
rect 4658 9222 4688 9274
rect 4688 9222 4700 9274
rect 4700 9222 4714 9274
rect 4738 9222 4752 9274
rect 4752 9222 4764 9274
rect 4764 9222 4794 9274
rect 4818 9222 4828 9274
rect 4828 9222 4874 9274
rect 4578 9220 4634 9222
rect 4658 9220 4714 9222
rect 4738 9220 4794 9222
rect 4818 9220 4874 9222
rect 5785 9818 5841 9820
rect 5865 9818 5921 9820
rect 5945 9818 6001 9820
rect 6025 9818 6081 9820
rect 5785 9766 5831 9818
rect 5831 9766 5841 9818
rect 5865 9766 5895 9818
rect 5895 9766 5907 9818
rect 5907 9766 5921 9818
rect 5945 9766 5959 9818
rect 5959 9766 5971 9818
rect 5971 9766 6001 9818
rect 6025 9766 6035 9818
rect 6035 9766 6081 9818
rect 5785 9764 5841 9766
rect 5865 9764 5921 9766
rect 5945 9764 6001 9766
rect 6025 9764 6081 9766
rect 6993 10362 7049 10364
rect 7073 10362 7129 10364
rect 7153 10362 7209 10364
rect 7233 10362 7289 10364
rect 6993 10310 7039 10362
rect 7039 10310 7049 10362
rect 7073 10310 7103 10362
rect 7103 10310 7115 10362
rect 7115 10310 7129 10362
rect 7153 10310 7167 10362
rect 7167 10310 7179 10362
rect 7179 10310 7209 10362
rect 7233 10310 7243 10362
rect 7243 10310 7289 10362
rect 6993 10308 7049 10310
rect 7073 10308 7129 10310
rect 7153 10308 7209 10310
rect 7233 10308 7289 10310
rect 3370 6554 3426 6556
rect 3450 6554 3506 6556
rect 3530 6554 3586 6556
rect 3610 6554 3666 6556
rect 3370 6502 3416 6554
rect 3416 6502 3426 6554
rect 3450 6502 3480 6554
rect 3480 6502 3492 6554
rect 3492 6502 3506 6554
rect 3530 6502 3544 6554
rect 3544 6502 3556 6554
rect 3556 6502 3586 6554
rect 3610 6502 3620 6554
rect 3620 6502 3666 6554
rect 3370 6500 3426 6502
rect 3450 6500 3506 6502
rect 3530 6500 3586 6502
rect 3610 6500 3666 6502
rect 4578 8186 4634 8188
rect 4658 8186 4714 8188
rect 4738 8186 4794 8188
rect 4818 8186 4874 8188
rect 4578 8134 4624 8186
rect 4624 8134 4634 8186
rect 4658 8134 4688 8186
rect 4688 8134 4700 8186
rect 4700 8134 4714 8186
rect 4738 8134 4752 8186
rect 4752 8134 4764 8186
rect 4764 8134 4794 8186
rect 4818 8134 4828 8186
rect 4828 8134 4874 8186
rect 4578 8132 4634 8134
rect 4658 8132 4714 8134
rect 4738 8132 4794 8134
rect 4818 8132 4874 8134
rect 5785 8730 5841 8732
rect 5865 8730 5921 8732
rect 5945 8730 6001 8732
rect 6025 8730 6081 8732
rect 5785 8678 5831 8730
rect 5831 8678 5841 8730
rect 5865 8678 5895 8730
rect 5895 8678 5907 8730
rect 5907 8678 5921 8730
rect 5945 8678 5959 8730
rect 5959 8678 5971 8730
rect 5971 8678 6001 8730
rect 6025 8678 6035 8730
rect 6035 8678 6081 8730
rect 5785 8676 5841 8678
rect 5865 8676 5921 8678
rect 5945 8676 6001 8678
rect 6025 8676 6081 8678
rect 6993 9274 7049 9276
rect 7073 9274 7129 9276
rect 7153 9274 7209 9276
rect 7233 9274 7289 9276
rect 6993 9222 7039 9274
rect 7039 9222 7049 9274
rect 7073 9222 7103 9274
rect 7103 9222 7115 9274
rect 7115 9222 7129 9274
rect 7153 9222 7167 9274
rect 7167 9222 7179 9274
rect 7179 9222 7209 9274
rect 7233 9222 7243 9274
rect 7243 9222 7289 9274
rect 6993 9220 7049 9222
rect 7073 9220 7129 9222
rect 7153 9220 7209 9222
rect 7233 9220 7289 9222
rect 5785 7642 5841 7644
rect 5865 7642 5921 7644
rect 5945 7642 6001 7644
rect 6025 7642 6081 7644
rect 5785 7590 5831 7642
rect 5831 7590 5841 7642
rect 5865 7590 5895 7642
rect 5895 7590 5907 7642
rect 5907 7590 5921 7642
rect 5945 7590 5959 7642
rect 5959 7590 5971 7642
rect 5971 7590 6001 7642
rect 6025 7590 6035 7642
rect 6035 7590 6081 7642
rect 5785 7588 5841 7590
rect 5865 7588 5921 7590
rect 5945 7588 6001 7590
rect 6025 7588 6081 7590
rect 4578 7098 4634 7100
rect 4658 7098 4714 7100
rect 4738 7098 4794 7100
rect 4818 7098 4874 7100
rect 4578 7046 4624 7098
rect 4624 7046 4634 7098
rect 4658 7046 4688 7098
rect 4688 7046 4700 7098
rect 4700 7046 4714 7098
rect 4738 7046 4752 7098
rect 4752 7046 4764 7098
rect 4764 7046 4794 7098
rect 4818 7046 4828 7098
rect 4828 7046 4874 7098
rect 4578 7044 4634 7046
rect 4658 7044 4714 7046
rect 4738 7044 4794 7046
rect 4818 7044 4874 7046
rect 3370 5466 3426 5468
rect 3450 5466 3506 5468
rect 3530 5466 3586 5468
rect 3610 5466 3666 5468
rect 3370 5414 3416 5466
rect 3416 5414 3426 5466
rect 3450 5414 3480 5466
rect 3480 5414 3492 5466
rect 3492 5414 3506 5466
rect 3530 5414 3544 5466
rect 3544 5414 3556 5466
rect 3556 5414 3586 5466
rect 3610 5414 3620 5466
rect 3620 5414 3666 5466
rect 3370 5412 3426 5414
rect 3450 5412 3506 5414
rect 3530 5412 3586 5414
rect 3610 5412 3666 5414
rect 3370 4378 3426 4380
rect 3450 4378 3506 4380
rect 3530 4378 3586 4380
rect 3610 4378 3666 4380
rect 3370 4326 3416 4378
rect 3416 4326 3426 4378
rect 3450 4326 3480 4378
rect 3480 4326 3492 4378
rect 3492 4326 3506 4378
rect 3530 4326 3544 4378
rect 3544 4326 3556 4378
rect 3556 4326 3586 4378
rect 3610 4326 3620 4378
rect 3620 4326 3666 4378
rect 3370 4324 3426 4326
rect 3450 4324 3506 4326
rect 3530 4324 3586 4326
rect 3610 4324 3666 4326
rect 3370 3290 3426 3292
rect 3450 3290 3506 3292
rect 3530 3290 3586 3292
rect 3610 3290 3666 3292
rect 3370 3238 3416 3290
rect 3416 3238 3426 3290
rect 3450 3238 3480 3290
rect 3480 3238 3492 3290
rect 3492 3238 3506 3290
rect 3530 3238 3544 3290
rect 3544 3238 3556 3290
rect 3556 3238 3586 3290
rect 3610 3238 3620 3290
rect 3620 3238 3666 3290
rect 3370 3236 3426 3238
rect 3450 3236 3506 3238
rect 3530 3236 3586 3238
rect 3610 3236 3666 3238
rect 2163 2746 2219 2748
rect 2243 2746 2299 2748
rect 2323 2746 2379 2748
rect 2403 2746 2459 2748
rect 2163 2694 2209 2746
rect 2209 2694 2219 2746
rect 2243 2694 2273 2746
rect 2273 2694 2285 2746
rect 2285 2694 2299 2746
rect 2323 2694 2337 2746
rect 2337 2694 2349 2746
rect 2349 2694 2379 2746
rect 2403 2694 2413 2746
rect 2413 2694 2459 2746
rect 2163 2692 2219 2694
rect 2243 2692 2299 2694
rect 2323 2692 2379 2694
rect 2403 2692 2459 2694
rect 4066 3440 4122 3496
rect 6993 8186 7049 8188
rect 7073 8186 7129 8188
rect 7153 8186 7209 8188
rect 7233 8186 7289 8188
rect 6993 8134 7039 8186
rect 7039 8134 7049 8186
rect 7073 8134 7103 8186
rect 7103 8134 7115 8186
rect 7115 8134 7129 8186
rect 7153 8134 7167 8186
rect 7167 8134 7179 8186
rect 7179 8134 7209 8186
rect 7233 8134 7243 8186
rect 7243 8134 7289 8186
rect 6993 8132 7049 8134
rect 7073 8132 7129 8134
rect 7153 8132 7209 8134
rect 7233 8132 7289 8134
rect 8200 10906 8256 10908
rect 8280 10906 8336 10908
rect 8360 10906 8416 10908
rect 8440 10906 8496 10908
rect 8200 10854 8246 10906
rect 8246 10854 8256 10906
rect 8280 10854 8310 10906
rect 8310 10854 8322 10906
rect 8322 10854 8336 10906
rect 8360 10854 8374 10906
rect 8374 10854 8386 10906
rect 8386 10854 8416 10906
rect 8440 10854 8450 10906
rect 8450 10854 8496 10906
rect 8200 10852 8256 10854
rect 8280 10852 8336 10854
rect 8360 10852 8416 10854
rect 8440 10852 8496 10854
rect 10615 10906 10671 10908
rect 10695 10906 10751 10908
rect 10775 10906 10831 10908
rect 10855 10906 10911 10908
rect 10615 10854 10661 10906
rect 10661 10854 10671 10906
rect 10695 10854 10725 10906
rect 10725 10854 10737 10906
rect 10737 10854 10751 10906
rect 10775 10854 10789 10906
rect 10789 10854 10801 10906
rect 10801 10854 10831 10906
rect 10855 10854 10865 10906
rect 10865 10854 10911 10906
rect 10615 10852 10671 10854
rect 10695 10852 10751 10854
rect 10775 10852 10831 10854
rect 10855 10852 10911 10854
rect 8200 9818 8256 9820
rect 8280 9818 8336 9820
rect 8360 9818 8416 9820
rect 8440 9818 8496 9820
rect 8200 9766 8246 9818
rect 8246 9766 8256 9818
rect 8280 9766 8310 9818
rect 8310 9766 8322 9818
rect 8322 9766 8336 9818
rect 8360 9766 8374 9818
rect 8374 9766 8386 9818
rect 8386 9766 8416 9818
rect 8440 9766 8450 9818
rect 8450 9766 8496 9818
rect 8200 9764 8256 9766
rect 8280 9764 8336 9766
rect 8360 9764 8416 9766
rect 8440 9764 8496 9766
rect 8200 8730 8256 8732
rect 8280 8730 8336 8732
rect 8360 8730 8416 8732
rect 8440 8730 8496 8732
rect 8200 8678 8246 8730
rect 8246 8678 8256 8730
rect 8280 8678 8310 8730
rect 8310 8678 8322 8730
rect 8322 8678 8336 8730
rect 8360 8678 8374 8730
rect 8374 8678 8386 8730
rect 8386 8678 8416 8730
rect 8440 8678 8450 8730
rect 8450 8678 8496 8730
rect 8200 8676 8256 8678
rect 8280 8676 8336 8678
rect 8360 8676 8416 8678
rect 8440 8676 8496 8678
rect 6993 7098 7049 7100
rect 7073 7098 7129 7100
rect 7153 7098 7209 7100
rect 7233 7098 7289 7100
rect 6993 7046 7039 7098
rect 7039 7046 7049 7098
rect 7073 7046 7103 7098
rect 7103 7046 7115 7098
rect 7115 7046 7129 7098
rect 7153 7046 7167 7098
rect 7167 7046 7179 7098
rect 7179 7046 7209 7098
rect 7233 7046 7243 7098
rect 7243 7046 7289 7098
rect 6993 7044 7049 7046
rect 7073 7044 7129 7046
rect 7153 7044 7209 7046
rect 7233 7044 7289 7046
rect 5785 6554 5841 6556
rect 5865 6554 5921 6556
rect 5945 6554 6001 6556
rect 6025 6554 6081 6556
rect 5785 6502 5831 6554
rect 5831 6502 5841 6554
rect 5865 6502 5895 6554
rect 5895 6502 5907 6554
rect 5907 6502 5921 6554
rect 5945 6502 5959 6554
rect 5959 6502 5971 6554
rect 5971 6502 6001 6554
rect 6025 6502 6035 6554
rect 6035 6502 6081 6554
rect 5785 6500 5841 6502
rect 5865 6500 5921 6502
rect 5945 6500 6001 6502
rect 6025 6500 6081 6502
rect 4578 6010 4634 6012
rect 4658 6010 4714 6012
rect 4738 6010 4794 6012
rect 4818 6010 4874 6012
rect 4578 5958 4624 6010
rect 4624 5958 4634 6010
rect 4658 5958 4688 6010
rect 4688 5958 4700 6010
rect 4700 5958 4714 6010
rect 4738 5958 4752 6010
rect 4752 5958 4764 6010
rect 4764 5958 4794 6010
rect 4818 5958 4828 6010
rect 4828 5958 4874 6010
rect 4578 5956 4634 5958
rect 4658 5956 4714 5958
rect 4738 5956 4794 5958
rect 4818 5956 4874 5958
rect 4578 4922 4634 4924
rect 4658 4922 4714 4924
rect 4738 4922 4794 4924
rect 4818 4922 4874 4924
rect 4578 4870 4624 4922
rect 4624 4870 4634 4922
rect 4658 4870 4688 4922
rect 4688 4870 4700 4922
rect 4700 4870 4714 4922
rect 4738 4870 4752 4922
rect 4752 4870 4764 4922
rect 4764 4870 4794 4922
rect 4818 4870 4828 4922
rect 4828 4870 4874 4922
rect 4578 4868 4634 4870
rect 4658 4868 4714 4870
rect 4738 4868 4794 4870
rect 4818 4868 4874 4870
rect 5785 5466 5841 5468
rect 5865 5466 5921 5468
rect 5945 5466 6001 5468
rect 6025 5466 6081 5468
rect 5785 5414 5831 5466
rect 5831 5414 5841 5466
rect 5865 5414 5895 5466
rect 5895 5414 5907 5466
rect 5907 5414 5921 5466
rect 5945 5414 5959 5466
rect 5959 5414 5971 5466
rect 5971 5414 6001 5466
rect 6025 5414 6035 5466
rect 6035 5414 6081 5466
rect 5785 5412 5841 5414
rect 5865 5412 5921 5414
rect 5945 5412 6001 5414
rect 6025 5412 6081 5414
rect 4578 3834 4634 3836
rect 4658 3834 4714 3836
rect 4738 3834 4794 3836
rect 4818 3834 4874 3836
rect 4578 3782 4624 3834
rect 4624 3782 4634 3834
rect 4658 3782 4688 3834
rect 4688 3782 4700 3834
rect 4700 3782 4714 3834
rect 4738 3782 4752 3834
rect 4752 3782 4764 3834
rect 4764 3782 4794 3834
rect 4818 3782 4828 3834
rect 4828 3782 4874 3834
rect 4578 3780 4634 3782
rect 4658 3780 4714 3782
rect 4738 3780 4794 3782
rect 4818 3780 4874 3782
rect 4578 2746 4634 2748
rect 4658 2746 4714 2748
rect 4738 2746 4794 2748
rect 4818 2746 4874 2748
rect 4578 2694 4624 2746
rect 4624 2694 4634 2746
rect 4658 2694 4688 2746
rect 4688 2694 4700 2746
rect 4700 2694 4714 2746
rect 4738 2694 4752 2746
rect 4752 2694 4764 2746
rect 4764 2694 4794 2746
rect 4818 2694 4828 2746
rect 4828 2694 4874 2746
rect 4578 2692 4634 2694
rect 4658 2692 4714 2694
rect 4738 2692 4794 2694
rect 4818 2692 4874 2694
rect 5785 4378 5841 4380
rect 5865 4378 5921 4380
rect 5945 4378 6001 4380
rect 6025 4378 6081 4380
rect 5785 4326 5831 4378
rect 5831 4326 5841 4378
rect 5865 4326 5895 4378
rect 5895 4326 5907 4378
rect 5907 4326 5921 4378
rect 5945 4326 5959 4378
rect 5959 4326 5971 4378
rect 5971 4326 6001 4378
rect 6025 4326 6035 4378
rect 6035 4326 6081 4378
rect 5785 4324 5841 4326
rect 5865 4324 5921 4326
rect 5945 4324 6001 4326
rect 6025 4324 6081 4326
rect 5785 3290 5841 3292
rect 5865 3290 5921 3292
rect 5945 3290 6001 3292
rect 6025 3290 6081 3292
rect 5785 3238 5831 3290
rect 5831 3238 5841 3290
rect 5865 3238 5895 3290
rect 5895 3238 5907 3290
rect 5907 3238 5921 3290
rect 5945 3238 5959 3290
rect 5959 3238 5971 3290
rect 5971 3238 6001 3290
rect 6025 3238 6035 3290
rect 6035 3238 6081 3290
rect 5785 3236 5841 3238
rect 5865 3236 5921 3238
rect 5945 3236 6001 3238
rect 6025 3236 6081 3238
rect 6993 6010 7049 6012
rect 7073 6010 7129 6012
rect 7153 6010 7209 6012
rect 7233 6010 7289 6012
rect 6993 5958 7039 6010
rect 7039 5958 7049 6010
rect 7073 5958 7103 6010
rect 7103 5958 7115 6010
rect 7115 5958 7129 6010
rect 7153 5958 7167 6010
rect 7167 5958 7179 6010
rect 7179 5958 7209 6010
rect 7233 5958 7243 6010
rect 7243 5958 7289 6010
rect 6993 5956 7049 5958
rect 7073 5956 7129 5958
rect 7153 5956 7209 5958
rect 7233 5956 7289 5958
rect 6993 4922 7049 4924
rect 7073 4922 7129 4924
rect 7153 4922 7209 4924
rect 7233 4922 7289 4924
rect 6993 4870 7039 4922
rect 7039 4870 7049 4922
rect 7073 4870 7103 4922
rect 7103 4870 7115 4922
rect 7115 4870 7129 4922
rect 7153 4870 7167 4922
rect 7167 4870 7179 4922
rect 7179 4870 7209 4922
rect 7233 4870 7243 4922
rect 7243 4870 7289 4922
rect 6993 4868 7049 4870
rect 7073 4868 7129 4870
rect 7153 4868 7209 4870
rect 7233 4868 7289 4870
rect 8200 7642 8256 7644
rect 8280 7642 8336 7644
rect 8360 7642 8416 7644
rect 8440 7642 8496 7644
rect 8200 7590 8246 7642
rect 8246 7590 8256 7642
rect 8280 7590 8310 7642
rect 8310 7590 8322 7642
rect 8322 7590 8336 7642
rect 8360 7590 8374 7642
rect 8374 7590 8386 7642
rect 8386 7590 8416 7642
rect 8440 7590 8450 7642
rect 8450 7590 8496 7642
rect 8200 7588 8256 7590
rect 8280 7588 8336 7590
rect 8360 7588 8416 7590
rect 8440 7588 8496 7590
rect 8200 6554 8256 6556
rect 8280 6554 8336 6556
rect 8360 6554 8416 6556
rect 8440 6554 8496 6556
rect 8200 6502 8246 6554
rect 8246 6502 8256 6554
rect 8280 6502 8310 6554
rect 8310 6502 8322 6554
rect 8322 6502 8336 6554
rect 8360 6502 8374 6554
rect 8374 6502 8386 6554
rect 8386 6502 8416 6554
rect 8440 6502 8450 6554
rect 8450 6502 8496 6554
rect 8200 6500 8256 6502
rect 8280 6500 8336 6502
rect 8360 6500 8416 6502
rect 8440 6500 8496 6502
rect 10874 10376 10930 10432
rect 9408 10362 9464 10364
rect 9488 10362 9544 10364
rect 9568 10362 9624 10364
rect 9648 10362 9704 10364
rect 9408 10310 9454 10362
rect 9454 10310 9464 10362
rect 9488 10310 9518 10362
rect 9518 10310 9530 10362
rect 9530 10310 9544 10362
rect 9568 10310 9582 10362
rect 9582 10310 9594 10362
rect 9594 10310 9624 10362
rect 9648 10310 9658 10362
rect 9658 10310 9704 10362
rect 9408 10308 9464 10310
rect 9488 10308 9544 10310
rect 9568 10308 9624 10310
rect 9648 10308 9704 10310
rect 9408 9274 9464 9276
rect 9488 9274 9544 9276
rect 9568 9274 9624 9276
rect 9648 9274 9704 9276
rect 9408 9222 9454 9274
rect 9454 9222 9464 9274
rect 9488 9222 9518 9274
rect 9518 9222 9530 9274
rect 9530 9222 9544 9274
rect 9568 9222 9582 9274
rect 9582 9222 9594 9274
rect 9594 9222 9624 9274
rect 9648 9222 9658 9274
rect 9658 9222 9704 9274
rect 9408 9220 9464 9222
rect 9488 9220 9544 9222
rect 9568 9220 9624 9222
rect 9648 9220 9704 9222
rect 9408 8186 9464 8188
rect 9488 8186 9544 8188
rect 9568 8186 9624 8188
rect 9648 8186 9704 8188
rect 9408 8134 9454 8186
rect 9454 8134 9464 8186
rect 9488 8134 9518 8186
rect 9518 8134 9530 8186
rect 9530 8134 9544 8186
rect 9568 8134 9582 8186
rect 9582 8134 9594 8186
rect 9594 8134 9624 8186
rect 9648 8134 9658 8186
rect 9658 8134 9704 8186
rect 9408 8132 9464 8134
rect 9488 8132 9544 8134
rect 9568 8132 9624 8134
rect 9648 8132 9704 8134
rect 9408 7098 9464 7100
rect 9488 7098 9544 7100
rect 9568 7098 9624 7100
rect 9648 7098 9704 7100
rect 9408 7046 9454 7098
rect 9454 7046 9464 7098
rect 9488 7046 9518 7098
rect 9518 7046 9530 7098
rect 9530 7046 9544 7098
rect 9568 7046 9582 7098
rect 9582 7046 9594 7098
rect 9594 7046 9624 7098
rect 9648 7046 9658 7098
rect 9658 7046 9704 7098
rect 9408 7044 9464 7046
rect 9488 7044 9544 7046
rect 9568 7044 9624 7046
rect 9648 7044 9704 7046
rect 6993 3834 7049 3836
rect 7073 3834 7129 3836
rect 7153 3834 7209 3836
rect 7233 3834 7289 3836
rect 6993 3782 7039 3834
rect 7039 3782 7049 3834
rect 7073 3782 7103 3834
rect 7103 3782 7115 3834
rect 7115 3782 7129 3834
rect 7153 3782 7167 3834
rect 7167 3782 7179 3834
rect 7179 3782 7209 3834
rect 7233 3782 7243 3834
rect 7243 3782 7289 3834
rect 6993 3780 7049 3782
rect 7073 3780 7129 3782
rect 7153 3780 7209 3782
rect 7233 3780 7289 3782
rect 8200 5466 8256 5468
rect 8280 5466 8336 5468
rect 8360 5466 8416 5468
rect 8440 5466 8496 5468
rect 8200 5414 8246 5466
rect 8246 5414 8256 5466
rect 8280 5414 8310 5466
rect 8310 5414 8322 5466
rect 8322 5414 8336 5466
rect 8360 5414 8374 5466
rect 8374 5414 8386 5466
rect 8386 5414 8416 5466
rect 8440 5414 8450 5466
rect 8450 5414 8496 5466
rect 8200 5412 8256 5414
rect 8280 5412 8336 5414
rect 8360 5412 8416 5414
rect 8440 5412 8496 5414
rect 8200 4378 8256 4380
rect 8280 4378 8336 4380
rect 8360 4378 8416 4380
rect 8440 4378 8496 4380
rect 8200 4326 8246 4378
rect 8246 4326 8256 4378
rect 8280 4326 8310 4378
rect 8310 4326 8322 4378
rect 8322 4326 8336 4378
rect 8360 4326 8374 4378
rect 8374 4326 8386 4378
rect 8386 4326 8416 4378
rect 8440 4326 8450 4378
rect 8450 4326 8496 4378
rect 8200 4324 8256 4326
rect 8280 4324 8336 4326
rect 8360 4324 8416 4326
rect 8440 4324 8496 4326
rect 6993 2746 7049 2748
rect 7073 2746 7129 2748
rect 7153 2746 7209 2748
rect 7233 2746 7289 2748
rect 6993 2694 7039 2746
rect 7039 2694 7049 2746
rect 7073 2694 7103 2746
rect 7103 2694 7115 2746
rect 7115 2694 7129 2746
rect 7153 2694 7167 2746
rect 7167 2694 7179 2746
rect 7179 2694 7209 2746
rect 7233 2694 7243 2746
rect 7243 2694 7289 2746
rect 6993 2692 7049 2694
rect 7073 2692 7129 2694
rect 7153 2692 7209 2694
rect 7233 2692 7289 2694
rect 8200 3290 8256 3292
rect 8280 3290 8336 3292
rect 8360 3290 8416 3292
rect 8440 3290 8496 3292
rect 8200 3238 8246 3290
rect 8246 3238 8256 3290
rect 8280 3238 8310 3290
rect 8310 3238 8322 3290
rect 8322 3238 8336 3290
rect 8360 3238 8374 3290
rect 8374 3238 8386 3290
rect 8386 3238 8416 3290
rect 8440 3238 8450 3290
rect 8450 3238 8496 3290
rect 8200 3236 8256 3238
rect 8280 3236 8336 3238
rect 8360 3236 8416 3238
rect 8440 3236 8496 3238
rect 3370 2202 3426 2204
rect 3450 2202 3506 2204
rect 3530 2202 3586 2204
rect 3610 2202 3666 2204
rect 3370 2150 3416 2202
rect 3416 2150 3426 2202
rect 3450 2150 3480 2202
rect 3480 2150 3492 2202
rect 3492 2150 3506 2202
rect 3530 2150 3544 2202
rect 3544 2150 3556 2202
rect 3556 2150 3586 2202
rect 3610 2150 3620 2202
rect 3620 2150 3666 2202
rect 3370 2148 3426 2150
rect 3450 2148 3506 2150
rect 3530 2148 3586 2150
rect 3610 2148 3666 2150
rect 5785 2202 5841 2204
rect 5865 2202 5921 2204
rect 5945 2202 6001 2204
rect 6025 2202 6081 2204
rect 5785 2150 5831 2202
rect 5831 2150 5841 2202
rect 5865 2150 5895 2202
rect 5895 2150 5907 2202
rect 5907 2150 5921 2202
rect 5945 2150 5959 2202
rect 5959 2150 5971 2202
rect 5971 2150 6001 2202
rect 6025 2150 6035 2202
rect 6035 2150 6081 2202
rect 5785 2148 5841 2150
rect 5865 2148 5921 2150
rect 5945 2148 6001 2150
rect 6025 2148 6081 2150
rect 8200 2202 8256 2204
rect 8280 2202 8336 2204
rect 8360 2202 8416 2204
rect 8440 2202 8496 2204
rect 8200 2150 8246 2202
rect 8246 2150 8256 2202
rect 8280 2150 8310 2202
rect 8310 2150 8322 2202
rect 8322 2150 8336 2202
rect 8360 2150 8374 2202
rect 8374 2150 8386 2202
rect 8386 2150 8416 2202
rect 8440 2150 8450 2202
rect 8450 2150 8496 2202
rect 8200 2148 8256 2150
rect 8280 2148 8336 2150
rect 8360 2148 8416 2150
rect 8440 2148 8496 2150
rect 9408 6010 9464 6012
rect 9488 6010 9544 6012
rect 9568 6010 9624 6012
rect 9648 6010 9704 6012
rect 9408 5958 9454 6010
rect 9454 5958 9464 6010
rect 9488 5958 9518 6010
rect 9518 5958 9530 6010
rect 9530 5958 9544 6010
rect 9568 5958 9582 6010
rect 9582 5958 9594 6010
rect 9594 5958 9624 6010
rect 9648 5958 9658 6010
rect 9658 5958 9704 6010
rect 9408 5956 9464 5958
rect 9488 5956 9544 5958
rect 9568 5956 9624 5958
rect 9648 5956 9704 5958
rect 9408 4922 9464 4924
rect 9488 4922 9544 4924
rect 9568 4922 9624 4924
rect 9648 4922 9704 4924
rect 9408 4870 9454 4922
rect 9454 4870 9464 4922
rect 9488 4870 9518 4922
rect 9518 4870 9530 4922
rect 9530 4870 9544 4922
rect 9568 4870 9582 4922
rect 9582 4870 9594 4922
rect 9594 4870 9624 4922
rect 9648 4870 9658 4922
rect 9658 4870 9704 4922
rect 9408 4868 9464 4870
rect 9488 4868 9544 4870
rect 9568 4868 9624 4870
rect 9648 4868 9704 4870
rect 9408 3834 9464 3836
rect 9488 3834 9544 3836
rect 9568 3834 9624 3836
rect 9648 3834 9704 3836
rect 9408 3782 9454 3834
rect 9454 3782 9464 3834
rect 9488 3782 9518 3834
rect 9518 3782 9530 3834
rect 9530 3782 9544 3834
rect 9568 3782 9582 3834
rect 9582 3782 9594 3834
rect 9594 3782 9624 3834
rect 9648 3782 9658 3834
rect 9658 3782 9704 3834
rect 9408 3780 9464 3782
rect 9488 3780 9544 3782
rect 9568 3780 9624 3782
rect 9648 3780 9704 3782
rect 9408 2746 9464 2748
rect 9488 2746 9544 2748
rect 9568 2746 9624 2748
rect 9648 2746 9704 2748
rect 9408 2694 9454 2746
rect 9454 2694 9464 2746
rect 9488 2694 9518 2746
rect 9518 2694 9530 2746
rect 9530 2694 9544 2746
rect 9568 2694 9582 2746
rect 9582 2694 9594 2746
rect 9594 2694 9624 2746
rect 9648 2694 9658 2746
rect 9658 2694 9704 2746
rect 9408 2692 9464 2694
rect 9488 2692 9544 2694
rect 9568 2692 9624 2694
rect 9648 2692 9704 2694
rect 10615 9818 10671 9820
rect 10695 9818 10751 9820
rect 10775 9818 10831 9820
rect 10855 9818 10911 9820
rect 10615 9766 10661 9818
rect 10661 9766 10671 9818
rect 10695 9766 10725 9818
rect 10725 9766 10737 9818
rect 10737 9766 10751 9818
rect 10775 9766 10789 9818
rect 10789 9766 10801 9818
rect 10801 9766 10831 9818
rect 10855 9766 10865 9818
rect 10865 9766 10911 9818
rect 10615 9764 10671 9766
rect 10695 9764 10751 9766
rect 10775 9764 10831 9766
rect 10855 9764 10911 9766
rect 10615 8730 10671 8732
rect 10695 8730 10751 8732
rect 10775 8730 10831 8732
rect 10855 8730 10911 8732
rect 10615 8678 10661 8730
rect 10661 8678 10671 8730
rect 10695 8678 10725 8730
rect 10725 8678 10737 8730
rect 10737 8678 10751 8730
rect 10775 8678 10789 8730
rect 10789 8678 10801 8730
rect 10801 8678 10831 8730
rect 10855 8678 10865 8730
rect 10865 8678 10911 8730
rect 10615 8676 10671 8678
rect 10695 8676 10751 8678
rect 10775 8676 10831 8678
rect 10855 8676 10911 8678
rect 10615 7642 10671 7644
rect 10695 7642 10751 7644
rect 10775 7642 10831 7644
rect 10855 7642 10911 7644
rect 10615 7590 10661 7642
rect 10661 7590 10671 7642
rect 10695 7590 10725 7642
rect 10725 7590 10737 7642
rect 10737 7590 10751 7642
rect 10775 7590 10789 7642
rect 10789 7590 10801 7642
rect 10801 7590 10831 7642
rect 10855 7590 10865 7642
rect 10865 7590 10911 7642
rect 10615 7588 10671 7590
rect 10695 7588 10751 7590
rect 10775 7588 10831 7590
rect 10855 7588 10911 7590
rect 10615 6554 10671 6556
rect 10695 6554 10751 6556
rect 10775 6554 10831 6556
rect 10855 6554 10911 6556
rect 10615 6502 10661 6554
rect 10661 6502 10671 6554
rect 10695 6502 10725 6554
rect 10725 6502 10737 6554
rect 10737 6502 10751 6554
rect 10775 6502 10789 6554
rect 10789 6502 10801 6554
rect 10801 6502 10831 6554
rect 10855 6502 10865 6554
rect 10865 6502 10911 6554
rect 10615 6500 10671 6502
rect 10695 6500 10751 6502
rect 10775 6500 10831 6502
rect 10855 6500 10911 6502
rect 10615 5466 10671 5468
rect 10695 5466 10751 5468
rect 10775 5466 10831 5468
rect 10855 5466 10911 5468
rect 10615 5414 10661 5466
rect 10661 5414 10671 5466
rect 10695 5414 10725 5466
rect 10725 5414 10737 5466
rect 10737 5414 10751 5466
rect 10775 5414 10789 5466
rect 10789 5414 10801 5466
rect 10801 5414 10831 5466
rect 10855 5414 10865 5466
rect 10865 5414 10911 5466
rect 10615 5412 10671 5414
rect 10695 5412 10751 5414
rect 10775 5412 10831 5414
rect 10855 5412 10911 5414
rect 10615 4378 10671 4380
rect 10695 4378 10751 4380
rect 10775 4378 10831 4380
rect 10855 4378 10911 4380
rect 10615 4326 10661 4378
rect 10661 4326 10671 4378
rect 10695 4326 10725 4378
rect 10725 4326 10737 4378
rect 10737 4326 10751 4378
rect 10775 4326 10789 4378
rect 10789 4326 10801 4378
rect 10801 4326 10831 4378
rect 10855 4326 10865 4378
rect 10865 4326 10911 4378
rect 10615 4324 10671 4326
rect 10695 4324 10751 4326
rect 10775 4324 10831 4326
rect 10855 4324 10911 4326
rect 10615 3290 10671 3292
rect 10695 3290 10751 3292
rect 10775 3290 10831 3292
rect 10855 3290 10911 3292
rect 10615 3238 10661 3290
rect 10661 3238 10671 3290
rect 10695 3238 10725 3290
rect 10725 3238 10737 3290
rect 10737 3238 10751 3290
rect 10775 3238 10789 3290
rect 10789 3238 10801 3290
rect 10801 3238 10831 3290
rect 10855 3238 10865 3290
rect 10865 3238 10911 3290
rect 10615 3236 10671 3238
rect 10695 3236 10751 3238
rect 10775 3236 10831 3238
rect 10855 3236 10911 3238
rect 10874 3052 10930 3088
rect 10874 3032 10876 3052
rect 10876 3032 10928 3052
rect 10928 3032 10930 3052
rect 10615 2202 10671 2204
rect 10695 2202 10751 2204
rect 10775 2202 10831 2204
rect 10855 2202 10911 2204
rect 10615 2150 10661 2202
rect 10661 2150 10671 2202
rect 10695 2150 10725 2202
rect 10725 2150 10737 2202
rect 10737 2150 10751 2202
rect 10775 2150 10789 2202
rect 10789 2150 10801 2202
rect 10801 2150 10831 2202
rect 10855 2150 10865 2202
rect 10865 2150 10911 2202
rect 10615 2148 10671 2150
rect 10695 2148 10751 2150
rect 10775 2148 10831 2150
rect 10855 2148 10911 2150
<< metal3 >>
rect 2153 11456 2469 11457
rect 2153 11392 2159 11456
rect 2223 11392 2239 11456
rect 2303 11392 2319 11456
rect 2383 11392 2399 11456
rect 2463 11392 2469 11456
rect 2153 11391 2469 11392
rect 4568 11456 4884 11457
rect 4568 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4814 11456
rect 4878 11392 4884 11456
rect 4568 11391 4884 11392
rect 6983 11456 7299 11457
rect 6983 11392 6989 11456
rect 7053 11392 7069 11456
rect 7133 11392 7149 11456
rect 7213 11392 7229 11456
rect 7293 11392 7299 11456
rect 6983 11391 7299 11392
rect 9398 11456 9714 11457
rect 9398 11392 9404 11456
rect 9468 11392 9484 11456
rect 9548 11392 9564 11456
rect 9628 11392 9644 11456
rect 9708 11392 9714 11456
rect 9398 11391 9714 11392
rect 3360 10912 3676 10913
rect 3360 10848 3366 10912
rect 3430 10848 3446 10912
rect 3510 10848 3526 10912
rect 3590 10848 3606 10912
rect 3670 10848 3676 10912
rect 3360 10847 3676 10848
rect 5775 10912 6091 10913
rect 5775 10848 5781 10912
rect 5845 10848 5861 10912
rect 5925 10848 5941 10912
rect 6005 10848 6021 10912
rect 6085 10848 6091 10912
rect 5775 10847 6091 10848
rect 8190 10912 8506 10913
rect 8190 10848 8196 10912
rect 8260 10848 8276 10912
rect 8340 10848 8356 10912
rect 8420 10848 8436 10912
rect 8500 10848 8506 10912
rect 8190 10847 8506 10848
rect 10605 10912 10921 10913
rect 10605 10848 10611 10912
rect 10675 10848 10691 10912
rect 10755 10848 10771 10912
rect 10835 10848 10851 10912
rect 10915 10848 10921 10912
rect 10605 10847 10921 10848
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 10869 10434 10935 10437
rect 11154 10434 11954 10464
rect 10869 10432 11954 10434
rect 10869 10376 10874 10432
rect 10930 10376 11954 10432
rect 10869 10374 11954 10376
rect 10869 10371 10935 10374
rect 2153 10368 2469 10369
rect 2153 10304 2159 10368
rect 2223 10304 2239 10368
rect 2303 10304 2319 10368
rect 2383 10304 2399 10368
rect 2463 10304 2469 10368
rect 2153 10303 2469 10304
rect 4568 10368 4884 10369
rect 4568 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4734 10368
rect 4798 10304 4814 10368
rect 4878 10304 4884 10368
rect 4568 10303 4884 10304
rect 6983 10368 7299 10369
rect 6983 10304 6989 10368
rect 7053 10304 7069 10368
rect 7133 10304 7149 10368
rect 7213 10304 7229 10368
rect 7293 10304 7299 10368
rect 6983 10303 7299 10304
rect 9398 10368 9714 10369
rect 9398 10304 9404 10368
rect 9468 10304 9484 10368
rect 9548 10304 9564 10368
rect 9628 10304 9644 10368
rect 9708 10304 9714 10368
rect 11154 10344 11954 10374
rect 9398 10303 9714 10304
rect 3360 9824 3676 9825
rect 3360 9760 3366 9824
rect 3430 9760 3446 9824
rect 3510 9760 3526 9824
rect 3590 9760 3606 9824
rect 3670 9760 3676 9824
rect 3360 9759 3676 9760
rect 5775 9824 6091 9825
rect 5775 9760 5781 9824
rect 5845 9760 5861 9824
rect 5925 9760 5941 9824
rect 6005 9760 6021 9824
rect 6085 9760 6091 9824
rect 5775 9759 6091 9760
rect 8190 9824 8506 9825
rect 8190 9760 8196 9824
rect 8260 9760 8276 9824
rect 8340 9760 8356 9824
rect 8420 9760 8436 9824
rect 8500 9760 8506 9824
rect 8190 9759 8506 9760
rect 10605 9824 10921 9825
rect 10605 9760 10611 9824
rect 10675 9760 10691 9824
rect 10755 9760 10771 9824
rect 10835 9760 10851 9824
rect 10915 9760 10921 9824
rect 10605 9759 10921 9760
rect 2153 9280 2469 9281
rect 2153 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2399 9280
rect 2463 9216 2469 9280
rect 2153 9215 2469 9216
rect 4568 9280 4884 9281
rect 4568 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4814 9280
rect 4878 9216 4884 9280
rect 4568 9215 4884 9216
rect 6983 9280 7299 9281
rect 6983 9216 6989 9280
rect 7053 9216 7069 9280
rect 7133 9216 7149 9280
rect 7213 9216 7229 9280
rect 7293 9216 7299 9280
rect 6983 9215 7299 9216
rect 9398 9280 9714 9281
rect 9398 9216 9404 9280
rect 9468 9216 9484 9280
rect 9548 9216 9564 9280
rect 9628 9216 9644 9280
rect 9708 9216 9714 9280
rect 9398 9215 9714 9216
rect 3360 8736 3676 8737
rect 3360 8672 3366 8736
rect 3430 8672 3446 8736
rect 3510 8672 3526 8736
rect 3590 8672 3606 8736
rect 3670 8672 3676 8736
rect 3360 8671 3676 8672
rect 5775 8736 6091 8737
rect 5775 8672 5781 8736
rect 5845 8672 5861 8736
rect 5925 8672 5941 8736
rect 6005 8672 6021 8736
rect 6085 8672 6091 8736
rect 5775 8671 6091 8672
rect 8190 8736 8506 8737
rect 8190 8672 8196 8736
rect 8260 8672 8276 8736
rect 8340 8672 8356 8736
rect 8420 8672 8436 8736
rect 8500 8672 8506 8736
rect 8190 8671 8506 8672
rect 10605 8736 10921 8737
rect 10605 8672 10611 8736
rect 10675 8672 10691 8736
rect 10755 8672 10771 8736
rect 10835 8672 10851 8736
rect 10915 8672 10921 8736
rect 10605 8671 10921 8672
rect 2153 8192 2469 8193
rect 2153 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2399 8192
rect 2463 8128 2469 8192
rect 2153 8127 2469 8128
rect 4568 8192 4884 8193
rect 4568 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4814 8192
rect 4878 8128 4884 8192
rect 4568 8127 4884 8128
rect 6983 8192 7299 8193
rect 6983 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7229 8192
rect 7293 8128 7299 8192
rect 6983 8127 7299 8128
rect 9398 8192 9714 8193
rect 9398 8128 9404 8192
rect 9468 8128 9484 8192
rect 9548 8128 9564 8192
rect 9628 8128 9644 8192
rect 9708 8128 9714 8192
rect 9398 8127 9714 8128
rect 3360 7648 3676 7649
rect 3360 7584 3366 7648
rect 3430 7584 3446 7648
rect 3510 7584 3526 7648
rect 3590 7584 3606 7648
rect 3670 7584 3676 7648
rect 3360 7583 3676 7584
rect 5775 7648 6091 7649
rect 5775 7584 5781 7648
rect 5845 7584 5861 7648
rect 5925 7584 5941 7648
rect 6005 7584 6021 7648
rect 6085 7584 6091 7648
rect 5775 7583 6091 7584
rect 8190 7648 8506 7649
rect 8190 7584 8196 7648
rect 8260 7584 8276 7648
rect 8340 7584 8356 7648
rect 8420 7584 8436 7648
rect 8500 7584 8506 7648
rect 8190 7583 8506 7584
rect 10605 7648 10921 7649
rect 10605 7584 10611 7648
rect 10675 7584 10691 7648
rect 10755 7584 10771 7648
rect 10835 7584 10851 7648
rect 10915 7584 10921 7648
rect 10605 7583 10921 7584
rect 2153 7104 2469 7105
rect 2153 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2399 7104
rect 2463 7040 2469 7104
rect 2153 7039 2469 7040
rect 4568 7104 4884 7105
rect 4568 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4814 7104
rect 4878 7040 4884 7104
rect 4568 7039 4884 7040
rect 6983 7104 7299 7105
rect 6983 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7229 7104
rect 7293 7040 7299 7104
rect 6983 7039 7299 7040
rect 9398 7104 9714 7105
rect 9398 7040 9404 7104
rect 9468 7040 9484 7104
rect 9548 7040 9564 7104
rect 9628 7040 9644 7104
rect 9708 7040 9714 7104
rect 9398 7039 9714 7040
rect 3360 6560 3676 6561
rect 3360 6496 3366 6560
rect 3430 6496 3446 6560
rect 3510 6496 3526 6560
rect 3590 6496 3606 6560
rect 3670 6496 3676 6560
rect 3360 6495 3676 6496
rect 5775 6560 6091 6561
rect 5775 6496 5781 6560
rect 5845 6496 5861 6560
rect 5925 6496 5941 6560
rect 6005 6496 6021 6560
rect 6085 6496 6091 6560
rect 5775 6495 6091 6496
rect 8190 6560 8506 6561
rect 8190 6496 8196 6560
rect 8260 6496 8276 6560
rect 8340 6496 8356 6560
rect 8420 6496 8436 6560
rect 8500 6496 8506 6560
rect 8190 6495 8506 6496
rect 10605 6560 10921 6561
rect 10605 6496 10611 6560
rect 10675 6496 10691 6560
rect 10755 6496 10771 6560
rect 10835 6496 10851 6560
rect 10915 6496 10921 6560
rect 10605 6495 10921 6496
rect 2153 6016 2469 6017
rect 2153 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2399 6016
rect 2463 5952 2469 6016
rect 2153 5951 2469 5952
rect 4568 6016 4884 6017
rect 4568 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4814 6016
rect 4878 5952 4884 6016
rect 4568 5951 4884 5952
rect 6983 6016 7299 6017
rect 6983 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7229 6016
rect 7293 5952 7299 6016
rect 6983 5951 7299 5952
rect 9398 6016 9714 6017
rect 9398 5952 9404 6016
rect 9468 5952 9484 6016
rect 9548 5952 9564 6016
rect 9628 5952 9644 6016
rect 9708 5952 9714 6016
rect 9398 5951 9714 5952
rect 3360 5472 3676 5473
rect 3360 5408 3366 5472
rect 3430 5408 3446 5472
rect 3510 5408 3526 5472
rect 3590 5408 3606 5472
rect 3670 5408 3676 5472
rect 3360 5407 3676 5408
rect 5775 5472 6091 5473
rect 5775 5408 5781 5472
rect 5845 5408 5861 5472
rect 5925 5408 5941 5472
rect 6005 5408 6021 5472
rect 6085 5408 6091 5472
rect 5775 5407 6091 5408
rect 8190 5472 8506 5473
rect 8190 5408 8196 5472
rect 8260 5408 8276 5472
rect 8340 5408 8356 5472
rect 8420 5408 8436 5472
rect 8500 5408 8506 5472
rect 8190 5407 8506 5408
rect 10605 5472 10921 5473
rect 10605 5408 10611 5472
rect 10675 5408 10691 5472
rect 10755 5408 10771 5472
rect 10835 5408 10851 5472
rect 10915 5408 10921 5472
rect 10605 5407 10921 5408
rect 2153 4928 2469 4929
rect 2153 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2399 4928
rect 2463 4864 2469 4928
rect 2153 4863 2469 4864
rect 4568 4928 4884 4929
rect 4568 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4814 4928
rect 4878 4864 4884 4928
rect 4568 4863 4884 4864
rect 6983 4928 7299 4929
rect 6983 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7229 4928
rect 7293 4864 7299 4928
rect 6983 4863 7299 4864
rect 9398 4928 9714 4929
rect 9398 4864 9404 4928
rect 9468 4864 9484 4928
rect 9548 4864 9564 4928
rect 9628 4864 9644 4928
rect 9708 4864 9714 4928
rect 9398 4863 9714 4864
rect 3360 4384 3676 4385
rect 3360 4320 3366 4384
rect 3430 4320 3446 4384
rect 3510 4320 3526 4384
rect 3590 4320 3606 4384
rect 3670 4320 3676 4384
rect 3360 4319 3676 4320
rect 5775 4384 6091 4385
rect 5775 4320 5781 4384
rect 5845 4320 5861 4384
rect 5925 4320 5941 4384
rect 6005 4320 6021 4384
rect 6085 4320 6091 4384
rect 5775 4319 6091 4320
rect 8190 4384 8506 4385
rect 8190 4320 8196 4384
rect 8260 4320 8276 4384
rect 8340 4320 8356 4384
rect 8420 4320 8436 4384
rect 8500 4320 8506 4384
rect 8190 4319 8506 4320
rect 10605 4384 10921 4385
rect 10605 4320 10611 4384
rect 10675 4320 10691 4384
rect 10755 4320 10771 4384
rect 10835 4320 10851 4384
rect 10915 4320 10921 4384
rect 10605 4319 10921 4320
rect 2153 3840 2469 3841
rect 2153 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2399 3840
rect 2463 3776 2469 3840
rect 2153 3775 2469 3776
rect 4568 3840 4884 3841
rect 4568 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4814 3840
rect 4878 3776 4884 3840
rect 4568 3775 4884 3776
rect 6983 3840 7299 3841
rect 6983 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7229 3840
rect 7293 3776 7299 3840
rect 6983 3775 7299 3776
rect 9398 3840 9714 3841
rect 9398 3776 9404 3840
rect 9468 3776 9484 3840
rect 9548 3776 9564 3840
rect 9628 3776 9644 3840
rect 9708 3776 9714 3840
rect 9398 3775 9714 3776
rect 4061 3498 4127 3501
rect 2638 3496 4127 3498
rect 2638 3440 4066 3496
rect 4122 3440 4127 3496
rect 2638 3438 4127 3440
rect 0 3362 800 3392
rect 2638 3362 2698 3438
rect 4061 3435 4127 3438
rect 11154 3362 11954 3392
rect 0 3302 2698 3362
rect 0 3272 800 3302
rect 3360 3296 3676 3297
rect 3360 3232 3366 3296
rect 3430 3232 3446 3296
rect 3510 3232 3526 3296
rect 3590 3232 3606 3296
rect 3670 3232 3676 3296
rect 3360 3231 3676 3232
rect 5775 3296 6091 3297
rect 5775 3232 5781 3296
rect 5845 3232 5861 3296
rect 5925 3232 5941 3296
rect 6005 3232 6021 3296
rect 6085 3232 6091 3296
rect 5775 3231 6091 3232
rect 8190 3296 8506 3297
rect 8190 3232 8196 3296
rect 8260 3232 8276 3296
rect 8340 3232 8356 3296
rect 8420 3232 8436 3296
rect 8500 3232 8506 3296
rect 8190 3231 8506 3232
rect 10605 3296 10921 3297
rect 10605 3232 10611 3296
rect 10675 3232 10691 3296
rect 10755 3232 10771 3296
rect 10835 3232 10851 3296
rect 10915 3232 10921 3296
rect 10605 3231 10921 3232
rect 11102 3272 11954 3362
rect 10869 3090 10935 3093
rect 11102 3090 11162 3272
rect 10869 3088 11162 3090
rect 10869 3032 10874 3088
rect 10930 3032 11162 3088
rect 10869 3030 11162 3032
rect 10869 3027 10935 3030
rect 2153 2752 2469 2753
rect 2153 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2399 2752
rect 2463 2688 2469 2752
rect 2153 2687 2469 2688
rect 4568 2752 4884 2753
rect 4568 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4814 2752
rect 4878 2688 4884 2752
rect 4568 2687 4884 2688
rect 6983 2752 7299 2753
rect 6983 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7229 2752
rect 7293 2688 7299 2752
rect 6983 2687 7299 2688
rect 9398 2752 9714 2753
rect 9398 2688 9404 2752
rect 9468 2688 9484 2752
rect 9548 2688 9564 2752
rect 9628 2688 9644 2752
rect 9708 2688 9714 2752
rect 9398 2687 9714 2688
rect 3360 2208 3676 2209
rect 3360 2144 3366 2208
rect 3430 2144 3446 2208
rect 3510 2144 3526 2208
rect 3590 2144 3606 2208
rect 3670 2144 3676 2208
rect 3360 2143 3676 2144
rect 5775 2208 6091 2209
rect 5775 2144 5781 2208
rect 5845 2144 5861 2208
rect 5925 2144 5941 2208
rect 6005 2144 6021 2208
rect 6085 2144 6091 2208
rect 5775 2143 6091 2144
rect 8190 2208 8506 2209
rect 8190 2144 8196 2208
rect 8260 2144 8276 2208
rect 8340 2144 8356 2208
rect 8420 2144 8436 2208
rect 8500 2144 8506 2208
rect 8190 2143 8506 2144
rect 10605 2208 10921 2209
rect 10605 2144 10611 2208
rect 10675 2144 10691 2208
rect 10755 2144 10771 2208
rect 10835 2144 10851 2208
rect 10915 2144 10921 2208
rect 10605 2143 10921 2144
<< via3 >>
rect 2159 11452 2223 11456
rect 2159 11396 2163 11452
rect 2163 11396 2219 11452
rect 2219 11396 2223 11452
rect 2159 11392 2223 11396
rect 2239 11452 2303 11456
rect 2239 11396 2243 11452
rect 2243 11396 2299 11452
rect 2299 11396 2303 11452
rect 2239 11392 2303 11396
rect 2319 11452 2383 11456
rect 2319 11396 2323 11452
rect 2323 11396 2379 11452
rect 2379 11396 2383 11452
rect 2319 11392 2383 11396
rect 2399 11452 2463 11456
rect 2399 11396 2403 11452
rect 2403 11396 2459 11452
rect 2459 11396 2463 11452
rect 2399 11392 2463 11396
rect 4574 11452 4638 11456
rect 4574 11396 4578 11452
rect 4578 11396 4634 11452
rect 4634 11396 4638 11452
rect 4574 11392 4638 11396
rect 4654 11452 4718 11456
rect 4654 11396 4658 11452
rect 4658 11396 4714 11452
rect 4714 11396 4718 11452
rect 4654 11392 4718 11396
rect 4734 11452 4798 11456
rect 4734 11396 4738 11452
rect 4738 11396 4794 11452
rect 4794 11396 4798 11452
rect 4734 11392 4798 11396
rect 4814 11452 4878 11456
rect 4814 11396 4818 11452
rect 4818 11396 4874 11452
rect 4874 11396 4878 11452
rect 4814 11392 4878 11396
rect 6989 11452 7053 11456
rect 6989 11396 6993 11452
rect 6993 11396 7049 11452
rect 7049 11396 7053 11452
rect 6989 11392 7053 11396
rect 7069 11452 7133 11456
rect 7069 11396 7073 11452
rect 7073 11396 7129 11452
rect 7129 11396 7133 11452
rect 7069 11392 7133 11396
rect 7149 11452 7213 11456
rect 7149 11396 7153 11452
rect 7153 11396 7209 11452
rect 7209 11396 7213 11452
rect 7149 11392 7213 11396
rect 7229 11452 7293 11456
rect 7229 11396 7233 11452
rect 7233 11396 7289 11452
rect 7289 11396 7293 11452
rect 7229 11392 7293 11396
rect 9404 11452 9468 11456
rect 9404 11396 9408 11452
rect 9408 11396 9464 11452
rect 9464 11396 9468 11452
rect 9404 11392 9468 11396
rect 9484 11452 9548 11456
rect 9484 11396 9488 11452
rect 9488 11396 9544 11452
rect 9544 11396 9548 11452
rect 9484 11392 9548 11396
rect 9564 11452 9628 11456
rect 9564 11396 9568 11452
rect 9568 11396 9624 11452
rect 9624 11396 9628 11452
rect 9564 11392 9628 11396
rect 9644 11452 9708 11456
rect 9644 11396 9648 11452
rect 9648 11396 9704 11452
rect 9704 11396 9708 11452
rect 9644 11392 9708 11396
rect 3366 10908 3430 10912
rect 3366 10852 3370 10908
rect 3370 10852 3426 10908
rect 3426 10852 3430 10908
rect 3366 10848 3430 10852
rect 3446 10908 3510 10912
rect 3446 10852 3450 10908
rect 3450 10852 3506 10908
rect 3506 10852 3510 10908
rect 3446 10848 3510 10852
rect 3526 10908 3590 10912
rect 3526 10852 3530 10908
rect 3530 10852 3586 10908
rect 3586 10852 3590 10908
rect 3526 10848 3590 10852
rect 3606 10908 3670 10912
rect 3606 10852 3610 10908
rect 3610 10852 3666 10908
rect 3666 10852 3670 10908
rect 3606 10848 3670 10852
rect 5781 10908 5845 10912
rect 5781 10852 5785 10908
rect 5785 10852 5841 10908
rect 5841 10852 5845 10908
rect 5781 10848 5845 10852
rect 5861 10908 5925 10912
rect 5861 10852 5865 10908
rect 5865 10852 5921 10908
rect 5921 10852 5925 10908
rect 5861 10848 5925 10852
rect 5941 10908 6005 10912
rect 5941 10852 5945 10908
rect 5945 10852 6001 10908
rect 6001 10852 6005 10908
rect 5941 10848 6005 10852
rect 6021 10908 6085 10912
rect 6021 10852 6025 10908
rect 6025 10852 6081 10908
rect 6081 10852 6085 10908
rect 6021 10848 6085 10852
rect 8196 10908 8260 10912
rect 8196 10852 8200 10908
rect 8200 10852 8256 10908
rect 8256 10852 8260 10908
rect 8196 10848 8260 10852
rect 8276 10908 8340 10912
rect 8276 10852 8280 10908
rect 8280 10852 8336 10908
rect 8336 10852 8340 10908
rect 8276 10848 8340 10852
rect 8356 10908 8420 10912
rect 8356 10852 8360 10908
rect 8360 10852 8416 10908
rect 8416 10852 8420 10908
rect 8356 10848 8420 10852
rect 8436 10908 8500 10912
rect 8436 10852 8440 10908
rect 8440 10852 8496 10908
rect 8496 10852 8500 10908
rect 8436 10848 8500 10852
rect 10611 10908 10675 10912
rect 10611 10852 10615 10908
rect 10615 10852 10671 10908
rect 10671 10852 10675 10908
rect 10611 10848 10675 10852
rect 10691 10908 10755 10912
rect 10691 10852 10695 10908
rect 10695 10852 10751 10908
rect 10751 10852 10755 10908
rect 10691 10848 10755 10852
rect 10771 10908 10835 10912
rect 10771 10852 10775 10908
rect 10775 10852 10831 10908
rect 10831 10852 10835 10908
rect 10771 10848 10835 10852
rect 10851 10908 10915 10912
rect 10851 10852 10855 10908
rect 10855 10852 10911 10908
rect 10911 10852 10915 10908
rect 10851 10848 10915 10852
rect 2159 10364 2223 10368
rect 2159 10308 2163 10364
rect 2163 10308 2219 10364
rect 2219 10308 2223 10364
rect 2159 10304 2223 10308
rect 2239 10364 2303 10368
rect 2239 10308 2243 10364
rect 2243 10308 2299 10364
rect 2299 10308 2303 10364
rect 2239 10304 2303 10308
rect 2319 10364 2383 10368
rect 2319 10308 2323 10364
rect 2323 10308 2379 10364
rect 2379 10308 2383 10364
rect 2319 10304 2383 10308
rect 2399 10364 2463 10368
rect 2399 10308 2403 10364
rect 2403 10308 2459 10364
rect 2459 10308 2463 10364
rect 2399 10304 2463 10308
rect 4574 10364 4638 10368
rect 4574 10308 4578 10364
rect 4578 10308 4634 10364
rect 4634 10308 4638 10364
rect 4574 10304 4638 10308
rect 4654 10364 4718 10368
rect 4654 10308 4658 10364
rect 4658 10308 4714 10364
rect 4714 10308 4718 10364
rect 4654 10304 4718 10308
rect 4734 10364 4798 10368
rect 4734 10308 4738 10364
rect 4738 10308 4794 10364
rect 4794 10308 4798 10364
rect 4734 10304 4798 10308
rect 4814 10364 4878 10368
rect 4814 10308 4818 10364
rect 4818 10308 4874 10364
rect 4874 10308 4878 10364
rect 4814 10304 4878 10308
rect 6989 10364 7053 10368
rect 6989 10308 6993 10364
rect 6993 10308 7049 10364
rect 7049 10308 7053 10364
rect 6989 10304 7053 10308
rect 7069 10364 7133 10368
rect 7069 10308 7073 10364
rect 7073 10308 7129 10364
rect 7129 10308 7133 10364
rect 7069 10304 7133 10308
rect 7149 10364 7213 10368
rect 7149 10308 7153 10364
rect 7153 10308 7209 10364
rect 7209 10308 7213 10364
rect 7149 10304 7213 10308
rect 7229 10364 7293 10368
rect 7229 10308 7233 10364
rect 7233 10308 7289 10364
rect 7289 10308 7293 10364
rect 7229 10304 7293 10308
rect 9404 10364 9468 10368
rect 9404 10308 9408 10364
rect 9408 10308 9464 10364
rect 9464 10308 9468 10364
rect 9404 10304 9468 10308
rect 9484 10364 9548 10368
rect 9484 10308 9488 10364
rect 9488 10308 9544 10364
rect 9544 10308 9548 10364
rect 9484 10304 9548 10308
rect 9564 10364 9628 10368
rect 9564 10308 9568 10364
rect 9568 10308 9624 10364
rect 9624 10308 9628 10364
rect 9564 10304 9628 10308
rect 9644 10364 9708 10368
rect 9644 10308 9648 10364
rect 9648 10308 9704 10364
rect 9704 10308 9708 10364
rect 9644 10304 9708 10308
rect 3366 9820 3430 9824
rect 3366 9764 3370 9820
rect 3370 9764 3426 9820
rect 3426 9764 3430 9820
rect 3366 9760 3430 9764
rect 3446 9820 3510 9824
rect 3446 9764 3450 9820
rect 3450 9764 3506 9820
rect 3506 9764 3510 9820
rect 3446 9760 3510 9764
rect 3526 9820 3590 9824
rect 3526 9764 3530 9820
rect 3530 9764 3586 9820
rect 3586 9764 3590 9820
rect 3526 9760 3590 9764
rect 3606 9820 3670 9824
rect 3606 9764 3610 9820
rect 3610 9764 3666 9820
rect 3666 9764 3670 9820
rect 3606 9760 3670 9764
rect 5781 9820 5845 9824
rect 5781 9764 5785 9820
rect 5785 9764 5841 9820
rect 5841 9764 5845 9820
rect 5781 9760 5845 9764
rect 5861 9820 5925 9824
rect 5861 9764 5865 9820
rect 5865 9764 5921 9820
rect 5921 9764 5925 9820
rect 5861 9760 5925 9764
rect 5941 9820 6005 9824
rect 5941 9764 5945 9820
rect 5945 9764 6001 9820
rect 6001 9764 6005 9820
rect 5941 9760 6005 9764
rect 6021 9820 6085 9824
rect 6021 9764 6025 9820
rect 6025 9764 6081 9820
rect 6081 9764 6085 9820
rect 6021 9760 6085 9764
rect 8196 9820 8260 9824
rect 8196 9764 8200 9820
rect 8200 9764 8256 9820
rect 8256 9764 8260 9820
rect 8196 9760 8260 9764
rect 8276 9820 8340 9824
rect 8276 9764 8280 9820
rect 8280 9764 8336 9820
rect 8336 9764 8340 9820
rect 8276 9760 8340 9764
rect 8356 9820 8420 9824
rect 8356 9764 8360 9820
rect 8360 9764 8416 9820
rect 8416 9764 8420 9820
rect 8356 9760 8420 9764
rect 8436 9820 8500 9824
rect 8436 9764 8440 9820
rect 8440 9764 8496 9820
rect 8496 9764 8500 9820
rect 8436 9760 8500 9764
rect 10611 9820 10675 9824
rect 10611 9764 10615 9820
rect 10615 9764 10671 9820
rect 10671 9764 10675 9820
rect 10611 9760 10675 9764
rect 10691 9820 10755 9824
rect 10691 9764 10695 9820
rect 10695 9764 10751 9820
rect 10751 9764 10755 9820
rect 10691 9760 10755 9764
rect 10771 9820 10835 9824
rect 10771 9764 10775 9820
rect 10775 9764 10831 9820
rect 10831 9764 10835 9820
rect 10771 9760 10835 9764
rect 10851 9820 10915 9824
rect 10851 9764 10855 9820
rect 10855 9764 10911 9820
rect 10911 9764 10915 9820
rect 10851 9760 10915 9764
rect 2159 9276 2223 9280
rect 2159 9220 2163 9276
rect 2163 9220 2219 9276
rect 2219 9220 2223 9276
rect 2159 9216 2223 9220
rect 2239 9276 2303 9280
rect 2239 9220 2243 9276
rect 2243 9220 2299 9276
rect 2299 9220 2303 9276
rect 2239 9216 2303 9220
rect 2319 9276 2383 9280
rect 2319 9220 2323 9276
rect 2323 9220 2379 9276
rect 2379 9220 2383 9276
rect 2319 9216 2383 9220
rect 2399 9276 2463 9280
rect 2399 9220 2403 9276
rect 2403 9220 2459 9276
rect 2459 9220 2463 9276
rect 2399 9216 2463 9220
rect 4574 9276 4638 9280
rect 4574 9220 4578 9276
rect 4578 9220 4634 9276
rect 4634 9220 4638 9276
rect 4574 9216 4638 9220
rect 4654 9276 4718 9280
rect 4654 9220 4658 9276
rect 4658 9220 4714 9276
rect 4714 9220 4718 9276
rect 4654 9216 4718 9220
rect 4734 9276 4798 9280
rect 4734 9220 4738 9276
rect 4738 9220 4794 9276
rect 4794 9220 4798 9276
rect 4734 9216 4798 9220
rect 4814 9276 4878 9280
rect 4814 9220 4818 9276
rect 4818 9220 4874 9276
rect 4874 9220 4878 9276
rect 4814 9216 4878 9220
rect 6989 9276 7053 9280
rect 6989 9220 6993 9276
rect 6993 9220 7049 9276
rect 7049 9220 7053 9276
rect 6989 9216 7053 9220
rect 7069 9276 7133 9280
rect 7069 9220 7073 9276
rect 7073 9220 7129 9276
rect 7129 9220 7133 9276
rect 7069 9216 7133 9220
rect 7149 9276 7213 9280
rect 7149 9220 7153 9276
rect 7153 9220 7209 9276
rect 7209 9220 7213 9276
rect 7149 9216 7213 9220
rect 7229 9276 7293 9280
rect 7229 9220 7233 9276
rect 7233 9220 7289 9276
rect 7289 9220 7293 9276
rect 7229 9216 7293 9220
rect 9404 9276 9468 9280
rect 9404 9220 9408 9276
rect 9408 9220 9464 9276
rect 9464 9220 9468 9276
rect 9404 9216 9468 9220
rect 9484 9276 9548 9280
rect 9484 9220 9488 9276
rect 9488 9220 9544 9276
rect 9544 9220 9548 9276
rect 9484 9216 9548 9220
rect 9564 9276 9628 9280
rect 9564 9220 9568 9276
rect 9568 9220 9624 9276
rect 9624 9220 9628 9276
rect 9564 9216 9628 9220
rect 9644 9276 9708 9280
rect 9644 9220 9648 9276
rect 9648 9220 9704 9276
rect 9704 9220 9708 9276
rect 9644 9216 9708 9220
rect 3366 8732 3430 8736
rect 3366 8676 3370 8732
rect 3370 8676 3426 8732
rect 3426 8676 3430 8732
rect 3366 8672 3430 8676
rect 3446 8732 3510 8736
rect 3446 8676 3450 8732
rect 3450 8676 3506 8732
rect 3506 8676 3510 8732
rect 3446 8672 3510 8676
rect 3526 8732 3590 8736
rect 3526 8676 3530 8732
rect 3530 8676 3586 8732
rect 3586 8676 3590 8732
rect 3526 8672 3590 8676
rect 3606 8732 3670 8736
rect 3606 8676 3610 8732
rect 3610 8676 3666 8732
rect 3666 8676 3670 8732
rect 3606 8672 3670 8676
rect 5781 8732 5845 8736
rect 5781 8676 5785 8732
rect 5785 8676 5841 8732
rect 5841 8676 5845 8732
rect 5781 8672 5845 8676
rect 5861 8732 5925 8736
rect 5861 8676 5865 8732
rect 5865 8676 5921 8732
rect 5921 8676 5925 8732
rect 5861 8672 5925 8676
rect 5941 8732 6005 8736
rect 5941 8676 5945 8732
rect 5945 8676 6001 8732
rect 6001 8676 6005 8732
rect 5941 8672 6005 8676
rect 6021 8732 6085 8736
rect 6021 8676 6025 8732
rect 6025 8676 6081 8732
rect 6081 8676 6085 8732
rect 6021 8672 6085 8676
rect 8196 8732 8260 8736
rect 8196 8676 8200 8732
rect 8200 8676 8256 8732
rect 8256 8676 8260 8732
rect 8196 8672 8260 8676
rect 8276 8732 8340 8736
rect 8276 8676 8280 8732
rect 8280 8676 8336 8732
rect 8336 8676 8340 8732
rect 8276 8672 8340 8676
rect 8356 8732 8420 8736
rect 8356 8676 8360 8732
rect 8360 8676 8416 8732
rect 8416 8676 8420 8732
rect 8356 8672 8420 8676
rect 8436 8732 8500 8736
rect 8436 8676 8440 8732
rect 8440 8676 8496 8732
rect 8496 8676 8500 8732
rect 8436 8672 8500 8676
rect 10611 8732 10675 8736
rect 10611 8676 10615 8732
rect 10615 8676 10671 8732
rect 10671 8676 10675 8732
rect 10611 8672 10675 8676
rect 10691 8732 10755 8736
rect 10691 8676 10695 8732
rect 10695 8676 10751 8732
rect 10751 8676 10755 8732
rect 10691 8672 10755 8676
rect 10771 8732 10835 8736
rect 10771 8676 10775 8732
rect 10775 8676 10831 8732
rect 10831 8676 10835 8732
rect 10771 8672 10835 8676
rect 10851 8732 10915 8736
rect 10851 8676 10855 8732
rect 10855 8676 10911 8732
rect 10911 8676 10915 8732
rect 10851 8672 10915 8676
rect 2159 8188 2223 8192
rect 2159 8132 2163 8188
rect 2163 8132 2219 8188
rect 2219 8132 2223 8188
rect 2159 8128 2223 8132
rect 2239 8188 2303 8192
rect 2239 8132 2243 8188
rect 2243 8132 2299 8188
rect 2299 8132 2303 8188
rect 2239 8128 2303 8132
rect 2319 8188 2383 8192
rect 2319 8132 2323 8188
rect 2323 8132 2379 8188
rect 2379 8132 2383 8188
rect 2319 8128 2383 8132
rect 2399 8188 2463 8192
rect 2399 8132 2403 8188
rect 2403 8132 2459 8188
rect 2459 8132 2463 8188
rect 2399 8128 2463 8132
rect 4574 8188 4638 8192
rect 4574 8132 4578 8188
rect 4578 8132 4634 8188
rect 4634 8132 4638 8188
rect 4574 8128 4638 8132
rect 4654 8188 4718 8192
rect 4654 8132 4658 8188
rect 4658 8132 4714 8188
rect 4714 8132 4718 8188
rect 4654 8128 4718 8132
rect 4734 8188 4798 8192
rect 4734 8132 4738 8188
rect 4738 8132 4794 8188
rect 4794 8132 4798 8188
rect 4734 8128 4798 8132
rect 4814 8188 4878 8192
rect 4814 8132 4818 8188
rect 4818 8132 4874 8188
rect 4874 8132 4878 8188
rect 4814 8128 4878 8132
rect 6989 8188 7053 8192
rect 6989 8132 6993 8188
rect 6993 8132 7049 8188
rect 7049 8132 7053 8188
rect 6989 8128 7053 8132
rect 7069 8188 7133 8192
rect 7069 8132 7073 8188
rect 7073 8132 7129 8188
rect 7129 8132 7133 8188
rect 7069 8128 7133 8132
rect 7149 8188 7213 8192
rect 7149 8132 7153 8188
rect 7153 8132 7209 8188
rect 7209 8132 7213 8188
rect 7149 8128 7213 8132
rect 7229 8188 7293 8192
rect 7229 8132 7233 8188
rect 7233 8132 7289 8188
rect 7289 8132 7293 8188
rect 7229 8128 7293 8132
rect 9404 8188 9468 8192
rect 9404 8132 9408 8188
rect 9408 8132 9464 8188
rect 9464 8132 9468 8188
rect 9404 8128 9468 8132
rect 9484 8188 9548 8192
rect 9484 8132 9488 8188
rect 9488 8132 9544 8188
rect 9544 8132 9548 8188
rect 9484 8128 9548 8132
rect 9564 8188 9628 8192
rect 9564 8132 9568 8188
rect 9568 8132 9624 8188
rect 9624 8132 9628 8188
rect 9564 8128 9628 8132
rect 9644 8188 9708 8192
rect 9644 8132 9648 8188
rect 9648 8132 9704 8188
rect 9704 8132 9708 8188
rect 9644 8128 9708 8132
rect 3366 7644 3430 7648
rect 3366 7588 3370 7644
rect 3370 7588 3426 7644
rect 3426 7588 3430 7644
rect 3366 7584 3430 7588
rect 3446 7644 3510 7648
rect 3446 7588 3450 7644
rect 3450 7588 3506 7644
rect 3506 7588 3510 7644
rect 3446 7584 3510 7588
rect 3526 7644 3590 7648
rect 3526 7588 3530 7644
rect 3530 7588 3586 7644
rect 3586 7588 3590 7644
rect 3526 7584 3590 7588
rect 3606 7644 3670 7648
rect 3606 7588 3610 7644
rect 3610 7588 3666 7644
rect 3666 7588 3670 7644
rect 3606 7584 3670 7588
rect 5781 7644 5845 7648
rect 5781 7588 5785 7644
rect 5785 7588 5841 7644
rect 5841 7588 5845 7644
rect 5781 7584 5845 7588
rect 5861 7644 5925 7648
rect 5861 7588 5865 7644
rect 5865 7588 5921 7644
rect 5921 7588 5925 7644
rect 5861 7584 5925 7588
rect 5941 7644 6005 7648
rect 5941 7588 5945 7644
rect 5945 7588 6001 7644
rect 6001 7588 6005 7644
rect 5941 7584 6005 7588
rect 6021 7644 6085 7648
rect 6021 7588 6025 7644
rect 6025 7588 6081 7644
rect 6081 7588 6085 7644
rect 6021 7584 6085 7588
rect 8196 7644 8260 7648
rect 8196 7588 8200 7644
rect 8200 7588 8256 7644
rect 8256 7588 8260 7644
rect 8196 7584 8260 7588
rect 8276 7644 8340 7648
rect 8276 7588 8280 7644
rect 8280 7588 8336 7644
rect 8336 7588 8340 7644
rect 8276 7584 8340 7588
rect 8356 7644 8420 7648
rect 8356 7588 8360 7644
rect 8360 7588 8416 7644
rect 8416 7588 8420 7644
rect 8356 7584 8420 7588
rect 8436 7644 8500 7648
rect 8436 7588 8440 7644
rect 8440 7588 8496 7644
rect 8496 7588 8500 7644
rect 8436 7584 8500 7588
rect 10611 7644 10675 7648
rect 10611 7588 10615 7644
rect 10615 7588 10671 7644
rect 10671 7588 10675 7644
rect 10611 7584 10675 7588
rect 10691 7644 10755 7648
rect 10691 7588 10695 7644
rect 10695 7588 10751 7644
rect 10751 7588 10755 7644
rect 10691 7584 10755 7588
rect 10771 7644 10835 7648
rect 10771 7588 10775 7644
rect 10775 7588 10831 7644
rect 10831 7588 10835 7644
rect 10771 7584 10835 7588
rect 10851 7644 10915 7648
rect 10851 7588 10855 7644
rect 10855 7588 10911 7644
rect 10911 7588 10915 7644
rect 10851 7584 10915 7588
rect 2159 7100 2223 7104
rect 2159 7044 2163 7100
rect 2163 7044 2219 7100
rect 2219 7044 2223 7100
rect 2159 7040 2223 7044
rect 2239 7100 2303 7104
rect 2239 7044 2243 7100
rect 2243 7044 2299 7100
rect 2299 7044 2303 7100
rect 2239 7040 2303 7044
rect 2319 7100 2383 7104
rect 2319 7044 2323 7100
rect 2323 7044 2379 7100
rect 2379 7044 2383 7100
rect 2319 7040 2383 7044
rect 2399 7100 2463 7104
rect 2399 7044 2403 7100
rect 2403 7044 2459 7100
rect 2459 7044 2463 7100
rect 2399 7040 2463 7044
rect 4574 7100 4638 7104
rect 4574 7044 4578 7100
rect 4578 7044 4634 7100
rect 4634 7044 4638 7100
rect 4574 7040 4638 7044
rect 4654 7100 4718 7104
rect 4654 7044 4658 7100
rect 4658 7044 4714 7100
rect 4714 7044 4718 7100
rect 4654 7040 4718 7044
rect 4734 7100 4798 7104
rect 4734 7044 4738 7100
rect 4738 7044 4794 7100
rect 4794 7044 4798 7100
rect 4734 7040 4798 7044
rect 4814 7100 4878 7104
rect 4814 7044 4818 7100
rect 4818 7044 4874 7100
rect 4874 7044 4878 7100
rect 4814 7040 4878 7044
rect 6989 7100 7053 7104
rect 6989 7044 6993 7100
rect 6993 7044 7049 7100
rect 7049 7044 7053 7100
rect 6989 7040 7053 7044
rect 7069 7100 7133 7104
rect 7069 7044 7073 7100
rect 7073 7044 7129 7100
rect 7129 7044 7133 7100
rect 7069 7040 7133 7044
rect 7149 7100 7213 7104
rect 7149 7044 7153 7100
rect 7153 7044 7209 7100
rect 7209 7044 7213 7100
rect 7149 7040 7213 7044
rect 7229 7100 7293 7104
rect 7229 7044 7233 7100
rect 7233 7044 7289 7100
rect 7289 7044 7293 7100
rect 7229 7040 7293 7044
rect 9404 7100 9468 7104
rect 9404 7044 9408 7100
rect 9408 7044 9464 7100
rect 9464 7044 9468 7100
rect 9404 7040 9468 7044
rect 9484 7100 9548 7104
rect 9484 7044 9488 7100
rect 9488 7044 9544 7100
rect 9544 7044 9548 7100
rect 9484 7040 9548 7044
rect 9564 7100 9628 7104
rect 9564 7044 9568 7100
rect 9568 7044 9624 7100
rect 9624 7044 9628 7100
rect 9564 7040 9628 7044
rect 9644 7100 9708 7104
rect 9644 7044 9648 7100
rect 9648 7044 9704 7100
rect 9704 7044 9708 7100
rect 9644 7040 9708 7044
rect 3366 6556 3430 6560
rect 3366 6500 3370 6556
rect 3370 6500 3426 6556
rect 3426 6500 3430 6556
rect 3366 6496 3430 6500
rect 3446 6556 3510 6560
rect 3446 6500 3450 6556
rect 3450 6500 3506 6556
rect 3506 6500 3510 6556
rect 3446 6496 3510 6500
rect 3526 6556 3590 6560
rect 3526 6500 3530 6556
rect 3530 6500 3586 6556
rect 3586 6500 3590 6556
rect 3526 6496 3590 6500
rect 3606 6556 3670 6560
rect 3606 6500 3610 6556
rect 3610 6500 3666 6556
rect 3666 6500 3670 6556
rect 3606 6496 3670 6500
rect 5781 6556 5845 6560
rect 5781 6500 5785 6556
rect 5785 6500 5841 6556
rect 5841 6500 5845 6556
rect 5781 6496 5845 6500
rect 5861 6556 5925 6560
rect 5861 6500 5865 6556
rect 5865 6500 5921 6556
rect 5921 6500 5925 6556
rect 5861 6496 5925 6500
rect 5941 6556 6005 6560
rect 5941 6500 5945 6556
rect 5945 6500 6001 6556
rect 6001 6500 6005 6556
rect 5941 6496 6005 6500
rect 6021 6556 6085 6560
rect 6021 6500 6025 6556
rect 6025 6500 6081 6556
rect 6081 6500 6085 6556
rect 6021 6496 6085 6500
rect 8196 6556 8260 6560
rect 8196 6500 8200 6556
rect 8200 6500 8256 6556
rect 8256 6500 8260 6556
rect 8196 6496 8260 6500
rect 8276 6556 8340 6560
rect 8276 6500 8280 6556
rect 8280 6500 8336 6556
rect 8336 6500 8340 6556
rect 8276 6496 8340 6500
rect 8356 6556 8420 6560
rect 8356 6500 8360 6556
rect 8360 6500 8416 6556
rect 8416 6500 8420 6556
rect 8356 6496 8420 6500
rect 8436 6556 8500 6560
rect 8436 6500 8440 6556
rect 8440 6500 8496 6556
rect 8496 6500 8500 6556
rect 8436 6496 8500 6500
rect 10611 6556 10675 6560
rect 10611 6500 10615 6556
rect 10615 6500 10671 6556
rect 10671 6500 10675 6556
rect 10611 6496 10675 6500
rect 10691 6556 10755 6560
rect 10691 6500 10695 6556
rect 10695 6500 10751 6556
rect 10751 6500 10755 6556
rect 10691 6496 10755 6500
rect 10771 6556 10835 6560
rect 10771 6500 10775 6556
rect 10775 6500 10831 6556
rect 10831 6500 10835 6556
rect 10771 6496 10835 6500
rect 10851 6556 10915 6560
rect 10851 6500 10855 6556
rect 10855 6500 10911 6556
rect 10911 6500 10915 6556
rect 10851 6496 10915 6500
rect 2159 6012 2223 6016
rect 2159 5956 2163 6012
rect 2163 5956 2219 6012
rect 2219 5956 2223 6012
rect 2159 5952 2223 5956
rect 2239 6012 2303 6016
rect 2239 5956 2243 6012
rect 2243 5956 2299 6012
rect 2299 5956 2303 6012
rect 2239 5952 2303 5956
rect 2319 6012 2383 6016
rect 2319 5956 2323 6012
rect 2323 5956 2379 6012
rect 2379 5956 2383 6012
rect 2319 5952 2383 5956
rect 2399 6012 2463 6016
rect 2399 5956 2403 6012
rect 2403 5956 2459 6012
rect 2459 5956 2463 6012
rect 2399 5952 2463 5956
rect 4574 6012 4638 6016
rect 4574 5956 4578 6012
rect 4578 5956 4634 6012
rect 4634 5956 4638 6012
rect 4574 5952 4638 5956
rect 4654 6012 4718 6016
rect 4654 5956 4658 6012
rect 4658 5956 4714 6012
rect 4714 5956 4718 6012
rect 4654 5952 4718 5956
rect 4734 6012 4798 6016
rect 4734 5956 4738 6012
rect 4738 5956 4794 6012
rect 4794 5956 4798 6012
rect 4734 5952 4798 5956
rect 4814 6012 4878 6016
rect 4814 5956 4818 6012
rect 4818 5956 4874 6012
rect 4874 5956 4878 6012
rect 4814 5952 4878 5956
rect 6989 6012 7053 6016
rect 6989 5956 6993 6012
rect 6993 5956 7049 6012
rect 7049 5956 7053 6012
rect 6989 5952 7053 5956
rect 7069 6012 7133 6016
rect 7069 5956 7073 6012
rect 7073 5956 7129 6012
rect 7129 5956 7133 6012
rect 7069 5952 7133 5956
rect 7149 6012 7213 6016
rect 7149 5956 7153 6012
rect 7153 5956 7209 6012
rect 7209 5956 7213 6012
rect 7149 5952 7213 5956
rect 7229 6012 7293 6016
rect 7229 5956 7233 6012
rect 7233 5956 7289 6012
rect 7289 5956 7293 6012
rect 7229 5952 7293 5956
rect 9404 6012 9468 6016
rect 9404 5956 9408 6012
rect 9408 5956 9464 6012
rect 9464 5956 9468 6012
rect 9404 5952 9468 5956
rect 9484 6012 9548 6016
rect 9484 5956 9488 6012
rect 9488 5956 9544 6012
rect 9544 5956 9548 6012
rect 9484 5952 9548 5956
rect 9564 6012 9628 6016
rect 9564 5956 9568 6012
rect 9568 5956 9624 6012
rect 9624 5956 9628 6012
rect 9564 5952 9628 5956
rect 9644 6012 9708 6016
rect 9644 5956 9648 6012
rect 9648 5956 9704 6012
rect 9704 5956 9708 6012
rect 9644 5952 9708 5956
rect 3366 5468 3430 5472
rect 3366 5412 3370 5468
rect 3370 5412 3426 5468
rect 3426 5412 3430 5468
rect 3366 5408 3430 5412
rect 3446 5468 3510 5472
rect 3446 5412 3450 5468
rect 3450 5412 3506 5468
rect 3506 5412 3510 5468
rect 3446 5408 3510 5412
rect 3526 5468 3590 5472
rect 3526 5412 3530 5468
rect 3530 5412 3586 5468
rect 3586 5412 3590 5468
rect 3526 5408 3590 5412
rect 3606 5468 3670 5472
rect 3606 5412 3610 5468
rect 3610 5412 3666 5468
rect 3666 5412 3670 5468
rect 3606 5408 3670 5412
rect 5781 5468 5845 5472
rect 5781 5412 5785 5468
rect 5785 5412 5841 5468
rect 5841 5412 5845 5468
rect 5781 5408 5845 5412
rect 5861 5468 5925 5472
rect 5861 5412 5865 5468
rect 5865 5412 5921 5468
rect 5921 5412 5925 5468
rect 5861 5408 5925 5412
rect 5941 5468 6005 5472
rect 5941 5412 5945 5468
rect 5945 5412 6001 5468
rect 6001 5412 6005 5468
rect 5941 5408 6005 5412
rect 6021 5468 6085 5472
rect 6021 5412 6025 5468
rect 6025 5412 6081 5468
rect 6081 5412 6085 5468
rect 6021 5408 6085 5412
rect 8196 5468 8260 5472
rect 8196 5412 8200 5468
rect 8200 5412 8256 5468
rect 8256 5412 8260 5468
rect 8196 5408 8260 5412
rect 8276 5468 8340 5472
rect 8276 5412 8280 5468
rect 8280 5412 8336 5468
rect 8336 5412 8340 5468
rect 8276 5408 8340 5412
rect 8356 5468 8420 5472
rect 8356 5412 8360 5468
rect 8360 5412 8416 5468
rect 8416 5412 8420 5468
rect 8356 5408 8420 5412
rect 8436 5468 8500 5472
rect 8436 5412 8440 5468
rect 8440 5412 8496 5468
rect 8496 5412 8500 5468
rect 8436 5408 8500 5412
rect 10611 5468 10675 5472
rect 10611 5412 10615 5468
rect 10615 5412 10671 5468
rect 10671 5412 10675 5468
rect 10611 5408 10675 5412
rect 10691 5468 10755 5472
rect 10691 5412 10695 5468
rect 10695 5412 10751 5468
rect 10751 5412 10755 5468
rect 10691 5408 10755 5412
rect 10771 5468 10835 5472
rect 10771 5412 10775 5468
rect 10775 5412 10831 5468
rect 10831 5412 10835 5468
rect 10771 5408 10835 5412
rect 10851 5468 10915 5472
rect 10851 5412 10855 5468
rect 10855 5412 10911 5468
rect 10911 5412 10915 5468
rect 10851 5408 10915 5412
rect 2159 4924 2223 4928
rect 2159 4868 2163 4924
rect 2163 4868 2219 4924
rect 2219 4868 2223 4924
rect 2159 4864 2223 4868
rect 2239 4924 2303 4928
rect 2239 4868 2243 4924
rect 2243 4868 2299 4924
rect 2299 4868 2303 4924
rect 2239 4864 2303 4868
rect 2319 4924 2383 4928
rect 2319 4868 2323 4924
rect 2323 4868 2379 4924
rect 2379 4868 2383 4924
rect 2319 4864 2383 4868
rect 2399 4924 2463 4928
rect 2399 4868 2403 4924
rect 2403 4868 2459 4924
rect 2459 4868 2463 4924
rect 2399 4864 2463 4868
rect 4574 4924 4638 4928
rect 4574 4868 4578 4924
rect 4578 4868 4634 4924
rect 4634 4868 4638 4924
rect 4574 4864 4638 4868
rect 4654 4924 4718 4928
rect 4654 4868 4658 4924
rect 4658 4868 4714 4924
rect 4714 4868 4718 4924
rect 4654 4864 4718 4868
rect 4734 4924 4798 4928
rect 4734 4868 4738 4924
rect 4738 4868 4794 4924
rect 4794 4868 4798 4924
rect 4734 4864 4798 4868
rect 4814 4924 4878 4928
rect 4814 4868 4818 4924
rect 4818 4868 4874 4924
rect 4874 4868 4878 4924
rect 4814 4864 4878 4868
rect 6989 4924 7053 4928
rect 6989 4868 6993 4924
rect 6993 4868 7049 4924
rect 7049 4868 7053 4924
rect 6989 4864 7053 4868
rect 7069 4924 7133 4928
rect 7069 4868 7073 4924
rect 7073 4868 7129 4924
rect 7129 4868 7133 4924
rect 7069 4864 7133 4868
rect 7149 4924 7213 4928
rect 7149 4868 7153 4924
rect 7153 4868 7209 4924
rect 7209 4868 7213 4924
rect 7149 4864 7213 4868
rect 7229 4924 7293 4928
rect 7229 4868 7233 4924
rect 7233 4868 7289 4924
rect 7289 4868 7293 4924
rect 7229 4864 7293 4868
rect 9404 4924 9468 4928
rect 9404 4868 9408 4924
rect 9408 4868 9464 4924
rect 9464 4868 9468 4924
rect 9404 4864 9468 4868
rect 9484 4924 9548 4928
rect 9484 4868 9488 4924
rect 9488 4868 9544 4924
rect 9544 4868 9548 4924
rect 9484 4864 9548 4868
rect 9564 4924 9628 4928
rect 9564 4868 9568 4924
rect 9568 4868 9624 4924
rect 9624 4868 9628 4924
rect 9564 4864 9628 4868
rect 9644 4924 9708 4928
rect 9644 4868 9648 4924
rect 9648 4868 9704 4924
rect 9704 4868 9708 4924
rect 9644 4864 9708 4868
rect 3366 4380 3430 4384
rect 3366 4324 3370 4380
rect 3370 4324 3426 4380
rect 3426 4324 3430 4380
rect 3366 4320 3430 4324
rect 3446 4380 3510 4384
rect 3446 4324 3450 4380
rect 3450 4324 3506 4380
rect 3506 4324 3510 4380
rect 3446 4320 3510 4324
rect 3526 4380 3590 4384
rect 3526 4324 3530 4380
rect 3530 4324 3586 4380
rect 3586 4324 3590 4380
rect 3526 4320 3590 4324
rect 3606 4380 3670 4384
rect 3606 4324 3610 4380
rect 3610 4324 3666 4380
rect 3666 4324 3670 4380
rect 3606 4320 3670 4324
rect 5781 4380 5845 4384
rect 5781 4324 5785 4380
rect 5785 4324 5841 4380
rect 5841 4324 5845 4380
rect 5781 4320 5845 4324
rect 5861 4380 5925 4384
rect 5861 4324 5865 4380
rect 5865 4324 5921 4380
rect 5921 4324 5925 4380
rect 5861 4320 5925 4324
rect 5941 4380 6005 4384
rect 5941 4324 5945 4380
rect 5945 4324 6001 4380
rect 6001 4324 6005 4380
rect 5941 4320 6005 4324
rect 6021 4380 6085 4384
rect 6021 4324 6025 4380
rect 6025 4324 6081 4380
rect 6081 4324 6085 4380
rect 6021 4320 6085 4324
rect 8196 4380 8260 4384
rect 8196 4324 8200 4380
rect 8200 4324 8256 4380
rect 8256 4324 8260 4380
rect 8196 4320 8260 4324
rect 8276 4380 8340 4384
rect 8276 4324 8280 4380
rect 8280 4324 8336 4380
rect 8336 4324 8340 4380
rect 8276 4320 8340 4324
rect 8356 4380 8420 4384
rect 8356 4324 8360 4380
rect 8360 4324 8416 4380
rect 8416 4324 8420 4380
rect 8356 4320 8420 4324
rect 8436 4380 8500 4384
rect 8436 4324 8440 4380
rect 8440 4324 8496 4380
rect 8496 4324 8500 4380
rect 8436 4320 8500 4324
rect 10611 4380 10675 4384
rect 10611 4324 10615 4380
rect 10615 4324 10671 4380
rect 10671 4324 10675 4380
rect 10611 4320 10675 4324
rect 10691 4380 10755 4384
rect 10691 4324 10695 4380
rect 10695 4324 10751 4380
rect 10751 4324 10755 4380
rect 10691 4320 10755 4324
rect 10771 4380 10835 4384
rect 10771 4324 10775 4380
rect 10775 4324 10831 4380
rect 10831 4324 10835 4380
rect 10771 4320 10835 4324
rect 10851 4380 10915 4384
rect 10851 4324 10855 4380
rect 10855 4324 10911 4380
rect 10911 4324 10915 4380
rect 10851 4320 10915 4324
rect 2159 3836 2223 3840
rect 2159 3780 2163 3836
rect 2163 3780 2219 3836
rect 2219 3780 2223 3836
rect 2159 3776 2223 3780
rect 2239 3836 2303 3840
rect 2239 3780 2243 3836
rect 2243 3780 2299 3836
rect 2299 3780 2303 3836
rect 2239 3776 2303 3780
rect 2319 3836 2383 3840
rect 2319 3780 2323 3836
rect 2323 3780 2379 3836
rect 2379 3780 2383 3836
rect 2319 3776 2383 3780
rect 2399 3836 2463 3840
rect 2399 3780 2403 3836
rect 2403 3780 2459 3836
rect 2459 3780 2463 3836
rect 2399 3776 2463 3780
rect 4574 3836 4638 3840
rect 4574 3780 4578 3836
rect 4578 3780 4634 3836
rect 4634 3780 4638 3836
rect 4574 3776 4638 3780
rect 4654 3836 4718 3840
rect 4654 3780 4658 3836
rect 4658 3780 4714 3836
rect 4714 3780 4718 3836
rect 4654 3776 4718 3780
rect 4734 3836 4798 3840
rect 4734 3780 4738 3836
rect 4738 3780 4794 3836
rect 4794 3780 4798 3836
rect 4734 3776 4798 3780
rect 4814 3836 4878 3840
rect 4814 3780 4818 3836
rect 4818 3780 4874 3836
rect 4874 3780 4878 3836
rect 4814 3776 4878 3780
rect 6989 3836 7053 3840
rect 6989 3780 6993 3836
rect 6993 3780 7049 3836
rect 7049 3780 7053 3836
rect 6989 3776 7053 3780
rect 7069 3836 7133 3840
rect 7069 3780 7073 3836
rect 7073 3780 7129 3836
rect 7129 3780 7133 3836
rect 7069 3776 7133 3780
rect 7149 3836 7213 3840
rect 7149 3780 7153 3836
rect 7153 3780 7209 3836
rect 7209 3780 7213 3836
rect 7149 3776 7213 3780
rect 7229 3836 7293 3840
rect 7229 3780 7233 3836
rect 7233 3780 7289 3836
rect 7289 3780 7293 3836
rect 7229 3776 7293 3780
rect 9404 3836 9468 3840
rect 9404 3780 9408 3836
rect 9408 3780 9464 3836
rect 9464 3780 9468 3836
rect 9404 3776 9468 3780
rect 9484 3836 9548 3840
rect 9484 3780 9488 3836
rect 9488 3780 9544 3836
rect 9544 3780 9548 3836
rect 9484 3776 9548 3780
rect 9564 3836 9628 3840
rect 9564 3780 9568 3836
rect 9568 3780 9624 3836
rect 9624 3780 9628 3836
rect 9564 3776 9628 3780
rect 9644 3836 9708 3840
rect 9644 3780 9648 3836
rect 9648 3780 9704 3836
rect 9704 3780 9708 3836
rect 9644 3776 9708 3780
rect 3366 3292 3430 3296
rect 3366 3236 3370 3292
rect 3370 3236 3426 3292
rect 3426 3236 3430 3292
rect 3366 3232 3430 3236
rect 3446 3292 3510 3296
rect 3446 3236 3450 3292
rect 3450 3236 3506 3292
rect 3506 3236 3510 3292
rect 3446 3232 3510 3236
rect 3526 3292 3590 3296
rect 3526 3236 3530 3292
rect 3530 3236 3586 3292
rect 3586 3236 3590 3292
rect 3526 3232 3590 3236
rect 3606 3292 3670 3296
rect 3606 3236 3610 3292
rect 3610 3236 3666 3292
rect 3666 3236 3670 3292
rect 3606 3232 3670 3236
rect 5781 3292 5845 3296
rect 5781 3236 5785 3292
rect 5785 3236 5841 3292
rect 5841 3236 5845 3292
rect 5781 3232 5845 3236
rect 5861 3292 5925 3296
rect 5861 3236 5865 3292
rect 5865 3236 5921 3292
rect 5921 3236 5925 3292
rect 5861 3232 5925 3236
rect 5941 3292 6005 3296
rect 5941 3236 5945 3292
rect 5945 3236 6001 3292
rect 6001 3236 6005 3292
rect 5941 3232 6005 3236
rect 6021 3292 6085 3296
rect 6021 3236 6025 3292
rect 6025 3236 6081 3292
rect 6081 3236 6085 3292
rect 6021 3232 6085 3236
rect 8196 3292 8260 3296
rect 8196 3236 8200 3292
rect 8200 3236 8256 3292
rect 8256 3236 8260 3292
rect 8196 3232 8260 3236
rect 8276 3292 8340 3296
rect 8276 3236 8280 3292
rect 8280 3236 8336 3292
rect 8336 3236 8340 3292
rect 8276 3232 8340 3236
rect 8356 3292 8420 3296
rect 8356 3236 8360 3292
rect 8360 3236 8416 3292
rect 8416 3236 8420 3292
rect 8356 3232 8420 3236
rect 8436 3292 8500 3296
rect 8436 3236 8440 3292
rect 8440 3236 8496 3292
rect 8496 3236 8500 3292
rect 8436 3232 8500 3236
rect 10611 3292 10675 3296
rect 10611 3236 10615 3292
rect 10615 3236 10671 3292
rect 10671 3236 10675 3292
rect 10611 3232 10675 3236
rect 10691 3292 10755 3296
rect 10691 3236 10695 3292
rect 10695 3236 10751 3292
rect 10751 3236 10755 3292
rect 10691 3232 10755 3236
rect 10771 3292 10835 3296
rect 10771 3236 10775 3292
rect 10775 3236 10831 3292
rect 10831 3236 10835 3292
rect 10771 3232 10835 3236
rect 10851 3292 10915 3296
rect 10851 3236 10855 3292
rect 10855 3236 10911 3292
rect 10911 3236 10915 3292
rect 10851 3232 10915 3236
rect 2159 2748 2223 2752
rect 2159 2692 2163 2748
rect 2163 2692 2219 2748
rect 2219 2692 2223 2748
rect 2159 2688 2223 2692
rect 2239 2748 2303 2752
rect 2239 2692 2243 2748
rect 2243 2692 2299 2748
rect 2299 2692 2303 2748
rect 2239 2688 2303 2692
rect 2319 2748 2383 2752
rect 2319 2692 2323 2748
rect 2323 2692 2379 2748
rect 2379 2692 2383 2748
rect 2319 2688 2383 2692
rect 2399 2748 2463 2752
rect 2399 2692 2403 2748
rect 2403 2692 2459 2748
rect 2459 2692 2463 2748
rect 2399 2688 2463 2692
rect 4574 2748 4638 2752
rect 4574 2692 4578 2748
rect 4578 2692 4634 2748
rect 4634 2692 4638 2748
rect 4574 2688 4638 2692
rect 4654 2748 4718 2752
rect 4654 2692 4658 2748
rect 4658 2692 4714 2748
rect 4714 2692 4718 2748
rect 4654 2688 4718 2692
rect 4734 2748 4798 2752
rect 4734 2692 4738 2748
rect 4738 2692 4794 2748
rect 4794 2692 4798 2748
rect 4734 2688 4798 2692
rect 4814 2748 4878 2752
rect 4814 2692 4818 2748
rect 4818 2692 4874 2748
rect 4874 2692 4878 2748
rect 4814 2688 4878 2692
rect 6989 2748 7053 2752
rect 6989 2692 6993 2748
rect 6993 2692 7049 2748
rect 7049 2692 7053 2748
rect 6989 2688 7053 2692
rect 7069 2748 7133 2752
rect 7069 2692 7073 2748
rect 7073 2692 7129 2748
rect 7129 2692 7133 2748
rect 7069 2688 7133 2692
rect 7149 2748 7213 2752
rect 7149 2692 7153 2748
rect 7153 2692 7209 2748
rect 7209 2692 7213 2748
rect 7149 2688 7213 2692
rect 7229 2748 7293 2752
rect 7229 2692 7233 2748
rect 7233 2692 7289 2748
rect 7289 2692 7293 2748
rect 7229 2688 7293 2692
rect 9404 2748 9468 2752
rect 9404 2692 9408 2748
rect 9408 2692 9464 2748
rect 9464 2692 9468 2748
rect 9404 2688 9468 2692
rect 9484 2748 9548 2752
rect 9484 2692 9488 2748
rect 9488 2692 9544 2748
rect 9544 2692 9548 2748
rect 9484 2688 9548 2692
rect 9564 2748 9628 2752
rect 9564 2692 9568 2748
rect 9568 2692 9624 2748
rect 9624 2692 9628 2748
rect 9564 2688 9628 2692
rect 9644 2748 9708 2752
rect 9644 2692 9648 2748
rect 9648 2692 9704 2748
rect 9704 2692 9708 2748
rect 9644 2688 9708 2692
rect 3366 2204 3430 2208
rect 3366 2148 3370 2204
rect 3370 2148 3426 2204
rect 3426 2148 3430 2204
rect 3366 2144 3430 2148
rect 3446 2204 3510 2208
rect 3446 2148 3450 2204
rect 3450 2148 3506 2204
rect 3506 2148 3510 2204
rect 3446 2144 3510 2148
rect 3526 2204 3590 2208
rect 3526 2148 3530 2204
rect 3530 2148 3586 2204
rect 3586 2148 3590 2204
rect 3526 2144 3590 2148
rect 3606 2204 3670 2208
rect 3606 2148 3610 2204
rect 3610 2148 3666 2204
rect 3666 2148 3670 2204
rect 3606 2144 3670 2148
rect 5781 2204 5845 2208
rect 5781 2148 5785 2204
rect 5785 2148 5841 2204
rect 5841 2148 5845 2204
rect 5781 2144 5845 2148
rect 5861 2204 5925 2208
rect 5861 2148 5865 2204
rect 5865 2148 5921 2204
rect 5921 2148 5925 2204
rect 5861 2144 5925 2148
rect 5941 2204 6005 2208
rect 5941 2148 5945 2204
rect 5945 2148 6001 2204
rect 6001 2148 6005 2204
rect 5941 2144 6005 2148
rect 6021 2204 6085 2208
rect 6021 2148 6025 2204
rect 6025 2148 6081 2204
rect 6081 2148 6085 2204
rect 6021 2144 6085 2148
rect 8196 2204 8260 2208
rect 8196 2148 8200 2204
rect 8200 2148 8256 2204
rect 8256 2148 8260 2204
rect 8196 2144 8260 2148
rect 8276 2204 8340 2208
rect 8276 2148 8280 2204
rect 8280 2148 8336 2204
rect 8336 2148 8340 2204
rect 8276 2144 8340 2148
rect 8356 2204 8420 2208
rect 8356 2148 8360 2204
rect 8360 2148 8416 2204
rect 8416 2148 8420 2204
rect 8356 2144 8420 2148
rect 8436 2204 8500 2208
rect 8436 2148 8440 2204
rect 8440 2148 8496 2204
rect 8496 2148 8500 2204
rect 8436 2144 8500 2148
rect 10611 2204 10675 2208
rect 10611 2148 10615 2204
rect 10615 2148 10671 2204
rect 10671 2148 10675 2204
rect 10611 2144 10675 2148
rect 10691 2204 10755 2208
rect 10691 2148 10695 2204
rect 10695 2148 10751 2204
rect 10751 2148 10755 2204
rect 10691 2144 10755 2148
rect 10771 2204 10835 2208
rect 10771 2148 10775 2204
rect 10775 2148 10831 2204
rect 10831 2148 10835 2204
rect 10771 2144 10835 2148
rect 10851 2204 10915 2208
rect 10851 2148 10855 2204
rect 10855 2148 10911 2204
rect 10911 2148 10915 2204
rect 10851 2144 10915 2148
<< metal4 >>
rect 2151 11456 2471 11472
rect 2151 11392 2159 11456
rect 2223 11392 2239 11456
rect 2303 11392 2319 11456
rect 2383 11392 2399 11456
rect 2463 11392 2471 11456
rect 2151 10368 2471 11392
rect 2151 10304 2159 10368
rect 2223 10304 2239 10368
rect 2303 10304 2319 10368
rect 2383 10304 2399 10368
rect 2463 10304 2471 10368
rect 2151 9280 2471 10304
rect 2151 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2399 9280
rect 2463 9216 2471 9280
rect 2151 8192 2471 9216
rect 2151 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2399 8192
rect 2463 8128 2471 8192
rect 2151 7104 2471 8128
rect 2151 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2399 7104
rect 2463 7040 2471 7104
rect 2151 6016 2471 7040
rect 2151 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2399 6016
rect 2463 5952 2471 6016
rect 2151 4928 2471 5952
rect 2151 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2399 4928
rect 2463 4864 2471 4928
rect 2151 3840 2471 4864
rect 2151 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2399 3840
rect 2463 3776 2471 3840
rect 2151 2752 2471 3776
rect 2151 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2399 2752
rect 2463 2688 2471 2752
rect 2151 2128 2471 2688
rect 3358 10912 3678 11472
rect 3358 10848 3366 10912
rect 3430 10848 3446 10912
rect 3510 10848 3526 10912
rect 3590 10848 3606 10912
rect 3670 10848 3678 10912
rect 3358 9824 3678 10848
rect 3358 9760 3366 9824
rect 3430 9760 3446 9824
rect 3510 9760 3526 9824
rect 3590 9760 3606 9824
rect 3670 9760 3678 9824
rect 3358 8736 3678 9760
rect 3358 8672 3366 8736
rect 3430 8672 3446 8736
rect 3510 8672 3526 8736
rect 3590 8672 3606 8736
rect 3670 8672 3678 8736
rect 3358 7648 3678 8672
rect 3358 7584 3366 7648
rect 3430 7584 3446 7648
rect 3510 7584 3526 7648
rect 3590 7584 3606 7648
rect 3670 7584 3678 7648
rect 3358 6560 3678 7584
rect 3358 6496 3366 6560
rect 3430 6496 3446 6560
rect 3510 6496 3526 6560
rect 3590 6496 3606 6560
rect 3670 6496 3678 6560
rect 3358 5472 3678 6496
rect 3358 5408 3366 5472
rect 3430 5408 3446 5472
rect 3510 5408 3526 5472
rect 3590 5408 3606 5472
rect 3670 5408 3678 5472
rect 3358 4384 3678 5408
rect 3358 4320 3366 4384
rect 3430 4320 3446 4384
rect 3510 4320 3526 4384
rect 3590 4320 3606 4384
rect 3670 4320 3678 4384
rect 3358 3296 3678 4320
rect 3358 3232 3366 3296
rect 3430 3232 3446 3296
rect 3510 3232 3526 3296
rect 3590 3232 3606 3296
rect 3670 3232 3678 3296
rect 3358 2208 3678 3232
rect 3358 2144 3366 2208
rect 3430 2144 3446 2208
rect 3510 2144 3526 2208
rect 3590 2144 3606 2208
rect 3670 2144 3678 2208
rect 3358 2128 3678 2144
rect 4566 11456 4886 11472
rect 4566 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4814 11456
rect 4878 11392 4886 11456
rect 4566 10368 4886 11392
rect 4566 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4734 10368
rect 4798 10304 4814 10368
rect 4878 10304 4886 10368
rect 4566 9280 4886 10304
rect 4566 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4814 9280
rect 4878 9216 4886 9280
rect 4566 8192 4886 9216
rect 4566 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4814 8192
rect 4878 8128 4886 8192
rect 4566 7104 4886 8128
rect 4566 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4814 7104
rect 4878 7040 4886 7104
rect 4566 6016 4886 7040
rect 4566 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4814 6016
rect 4878 5952 4886 6016
rect 4566 4928 4886 5952
rect 4566 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4814 4928
rect 4878 4864 4886 4928
rect 4566 3840 4886 4864
rect 4566 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4814 3840
rect 4878 3776 4886 3840
rect 4566 2752 4886 3776
rect 4566 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4814 2752
rect 4878 2688 4886 2752
rect 4566 2128 4886 2688
rect 5773 10912 6093 11472
rect 5773 10848 5781 10912
rect 5845 10848 5861 10912
rect 5925 10848 5941 10912
rect 6005 10848 6021 10912
rect 6085 10848 6093 10912
rect 5773 9824 6093 10848
rect 5773 9760 5781 9824
rect 5845 9760 5861 9824
rect 5925 9760 5941 9824
rect 6005 9760 6021 9824
rect 6085 9760 6093 9824
rect 5773 8736 6093 9760
rect 5773 8672 5781 8736
rect 5845 8672 5861 8736
rect 5925 8672 5941 8736
rect 6005 8672 6021 8736
rect 6085 8672 6093 8736
rect 5773 7648 6093 8672
rect 5773 7584 5781 7648
rect 5845 7584 5861 7648
rect 5925 7584 5941 7648
rect 6005 7584 6021 7648
rect 6085 7584 6093 7648
rect 5773 6560 6093 7584
rect 5773 6496 5781 6560
rect 5845 6496 5861 6560
rect 5925 6496 5941 6560
rect 6005 6496 6021 6560
rect 6085 6496 6093 6560
rect 5773 5472 6093 6496
rect 5773 5408 5781 5472
rect 5845 5408 5861 5472
rect 5925 5408 5941 5472
rect 6005 5408 6021 5472
rect 6085 5408 6093 5472
rect 5773 4384 6093 5408
rect 5773 4320 5781 4384
rect 5845 4320 5861 4384
rect 5925 4320 5941 4384
rect 6005 4320 6021 4384
rect 6085 4320 6093 4384
rect 5773 3296 6093 4320
rect 5773 3232 5781 3296
rect 5845 3232 5861 3296
rect 5925 3232 5941 3296
rect 6005 3232 6021 3296
rect 6085 3232 6093 3296
rect 5773 2208 6093 3232
rect 5773 2144 5781 2208
rect 5845 2144 5861 2208
rect 5925 2144 5941 2208
rect 6005 2144 6021 2208
rect 6085 2144 6093 2208
rect 5773 2128 6093 2144
rect 6981 11456 7301 11472
rect 6981 11392 6989 11456
rect 7053 11392 7069 11456
rect 7133 11392 7149 11456
rect 7213 11392 7229 11456
rect 7293 11392 7301 11456
rect 6981 10368 7301 11392
rect 6981 10304 6989 10368
rect 7053 10304 7069 10368
rect 7133 10304 7149 10368
rect 7213 10304 7229 10368
rect 7293 10304 7301 10368
rect 6981 9280 7301 10304
rect 6981 9216 6989 9280
rect 7053 9216 7069 9280
rect 7133 9216 7149 9280
rect 7213 9216 7229 9280
rect 7293 9216 7301 9280
rect 6981 8192 7301 9216
rect 6981 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7229 8192
rect 7293 8128 7301 8192
rect 6981 7104 7301 8128
rect 6981 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7229 7104
rect 7293 7040 7301 7104
rect 6981 6016 7301 7040
rect 6981 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7229 6016
rect 7293 5952 7301 6016
rect 6981 4928 7301 5952
rect 6981 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7229 4928
rect 7293 4864 7301 4928
rect 6981 3840 7301 4864
rect 6981 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7229 3840
rect 7293 3776 7301 3840
rect 6981 2752 7301 3776
rect 6981 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7229 2752
rect 7293 2688 7301 2752
rect 6981 2128 7301 2688
rect 8188 10912 8508 11472
rect 8188 10848 8196 10912
rect 8260 10848 8276 10912
rect 8340 10848 8356 10912
rect 8420 10848 8436 10912
rect 8500 10848 8508 10912
rect 8188 9824 8508 10848
rect 8188 9760 8196 9824
rect 8260 9760 8276 9824
rect 8340 9760 8356 9824
rect 8420 9760 8436 9824
rect 8500 9760 8508 9824
rect 8188 8736 8508 9760
rect 8188 8672 8196 8736
rect 8260 8672 8276 8736
rect 8340 8672 8356 8736
rect 8420 8672 8436 8736
rect 8500 8672 8508 8736
rect 8188 7648 8508 8672
rect 8188 7584 8196 7648
rect 8260 7584 8276 7648
rect 8340 7584 8356 7648
rect 8420 7584 8436 7648
rect 8500 7584 8508 7648
rect 8188 6560 8508 7584
rect 8188 6496 8196 6560
rect 8260 6496 8276 6560
rect 8340 6496 8356 6560
rect 8420 6496 8436 6560
rect 8500 6496 8508 6560
rect 8188 5472 8508 6496
rect 8188 5408 8196 5472
rect 8260 5408 8276 5472
rect 8340 5408 8356 5472
rect 8420 5408 8436 5472
rect 8500 5408 8508 5472
rect 8188 4384 8508 5408
rect 8188 4320 8196 4384
rect 8260 4320 8276 4384
rect 8340 4320 8356 4384
rect 8420 4320 8436 4384
rect 8500 4320 8508 4384
rect 8188 3296 8508 4320
rect 8188 3232 8196 3296
rect 8260 3232 8276 3296
rect 8340 3232 8356 3296
rect 8420 3232 8436 3296
rect 8500 3232 8508 3296
rect 8188 2208 8508 3232
rect 8188 2144 8196 2208
rect 8260 2144 8276 2208
rect 8340 2144 8356 2208
rect 8420 2144 8436 2208
rect 8500 2144 8508 2208
rect 8188 2128 8508 2144
rect 9396 11456 9716 11472
rect 9396 11392 9404 11456
rect 9468 11392 9484 11456
rect 9548 11392 9564 11456
rect 9628 11392 9644 11456
rect 9708 11392 9716 11456
rect 9396 10368 9716 11392
rect 9396 10304 9404 10368
rect 9468 10304 9484 10368
rect 9548 10304 9564 10368
rect 9628 10304 9644 10368
rect 9708 10304 9716 10368
rect 9396 9280 9716 10304
rect 9396 9216 9404 9280
rect 9468 9216 9484 9280
rect 9548 9216 9564 9280
rect 9628 9216 9644 9280
rect 9708 9216 9716 9280
rect 9396 8192 9716 9216
rect 9396 8128 9404 8192
rect 9468 8128 9484 8192
rect 9548 8128 9564 8192
rect 9628 8128 9644 8192
rect 9708 8128 9716 8192
rect 9396 7104 9716 8128
rect 9396 7040 9404 7104
rect 9468 7040 9484 7104
rect 9548 7040 9564 7104
rect 9628 7040 9644 7104
rect 9708 7040 9716 7104
rect 9396 6016 9716 7040
rect 9396 5952 9404 6016
rect 9468 5952 9484 6016
rect 9548 5952 9564 6016
rect 9628 5952 9644 6016
rect 9708 5952 9716 6016
rect 9396 4928 9716 5952
rect 9396 4864 9404 4928
rect 9468 4864 9484 4928
rect 9548 4864 9564 4928
rect 9628 4864 9644 4928
rect 9708 4864 9716 4928
rect 9396 3840 9716 4864
rect 9396 3776 9404 3840
rect 9468 3776 9484 3840
rect 9548 3776 9564 3840
rect 9628 3776 9644 3840
rect 9708 3776 9716 3840
rect 9396 2752 9716 3776
rect 9396 2688 9404 2752
rect 9468 2688 9484 2752
rect 9548 2688 9564 2752
rect 9628 2688 9644 2752
rect 9708 2688 9716 2752
rect 9396 2128 9716 2688
rect 10603 10912 10923 11472
rect 10603 10848 10611 10912
rect 10675 10848 10691 10912
rect 10755 10848 10771 10912
rect 10835 10848 10851 10912
rect 10915 10848 10923 10912
rect 10603 9824 10923 10848
rect 10603 9760 10611 9824
rect 10675 9760 10691 9824
rect 10755 9760 10771 9824
rect 10835 9760 10851 9824
rect 10915 9760 10923 9824
rect 10603 8736 10923 9760
rect 10603 8672 10611 8736
rect 10675 8672 10691 8736
rect 10755 8672 10771 8736
rect 10835 8672 10851 8736
rect 10915 8672 10923 8736
rect 10603 7648 10923 8672
rect 10603 7584 10611 7648
rect 10675 7584 10691 7648
rect 10755 7584 10771 7648
rect 10835 7584 10851 7648
rect 10915 7584 10923 7648
rect 10603 6560 10923 7584
rect 10603 6496 10611 6560
rect 10675 6496 10691 6560
rect 10755 6496 10771 6560
rect 10835 6496 10851 6560
rect 10915 6496 10923 6560
rect 10603 5472 10923 6496
rect 10603 5408 10611 5472
rect 10675 5408 10691 5472
rect 10755 5408 10771 5472
rect 10835 5408 10851 5472
rect 10915 5408 10923 5472
rect 10603 4384 10923 5408
rect 10603 4320 10611 4384
rect 10675 4320 10691 4384
rect 10755 4320 10771 4384
rect 10835 4320 10851 4384
rect 10915 4320 10923 4384
rect 10603 3296 10923 4320
rect 10603 3232 10611 3296
rect 10675 3232 10691 3296
rect 10755 3232 10771 3296
rect 10835 3232 10851 3296
rect 10915 3232 10923 3296
rect 10603 2208 10923 3232
rect 10603 2144 10611 2208
rect 10675 2144 10691 2208
rect 10755 2144 10771 2208
rect 10835 2144 10851 2208
rect 10915 2144 10923 2208
rect 10603 2128 10923 2144
use sky130_fd_sc_hd__or3b_1  _049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 4232 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 5152 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5980 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _053_
timestamp 1717180972
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1717180972
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1717180972
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 4416 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _058_
timestamp 1717180972
transform 1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _059_
timestamp 1717180972
transform 1 0 3772 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _060_
timestamp 1717180972
transform -1 0 3772 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _063_
timestamp 1717180972
transform -1 0 10396 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _065_
timestamp 1717180972
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10028 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 8096 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _071_
timestamp 1717180972
transform -1 0 8740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 7636 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1717180972
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _074_
timestamp 1717180972
transform 1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _075_
timestamp 1717180972
transform 1 0 8004 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _076_
timestamp 1717180972
transform 1 0 3128 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _077_
timestamp 1717180972
transform -1 0 4416 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _078_
timestamp 1717180972
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _079_
timestamp 1717180972
transform -1 0 3680 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _080_
timestamp 1717180972
transform -1 0 2208 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _082_
timestamp 1717180972
transform -1 0 2392 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _083_
timestamp 1717180972
transform -1 0 2484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1717180972
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 9936 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _087_
timestamp 1717180972
transform 1 0 8372 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _088_
timestamp 1717180972
transform -1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _089_
timestamp 1717180972
transform -1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1717180972
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1717180972
transform -1 0 8740 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1717180972
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _093_
timestamp 1717180972
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _095_
timestamp 1717180972
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _096_
timestamp 1717180972
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7268 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 6072 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _099_
timestamp 1717180972
transform 1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _103_
timestamp 1717180972
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp 1717180972
transform 1 0 8464 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp 1717180972
transform 1 0 9016 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _107_
timestamp 1717180972
transform 1 0 7084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 1717180972
transform 1 0 7636 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _109_
timestamp 1717180972
transform 1 0 3772 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _110_
timestamp 1717180972
transform 1 0 1932 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _111_
timestamp 1717180972
transform -1 0 5796 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp 1717180972
transform 1 0 3772 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp 1717180972
transform 1 0 1564 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp 1717180972
transform 1 0 1656 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _115_
timestamp 1717180972
transform 1 0 9016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _116_
timestamp 1717180972
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 1717180972
transform 1 0 5244 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 1717180972
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp 1717180972
transform 1 0 5520 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _120_
timestamp 1717180972
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 1717180972
transform -1 0 5704 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 1717180972
transform 1 0 6256 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _123_
timestamp 1717180972
transform 1 0 9016 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 1717180972
transform 1 0 7912 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 5336 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1717180972
transform -1 0 6256 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1717180972
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 1717180972
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1717180972
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1717180972
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_11
timestamp 1717180972
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_29
timestamp 1717180972
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1717180972
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1717180972
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1717180972
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1717180972
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_96
timestamp 1717180972
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1717180972
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1717180972
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1717180972
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1717180972
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 1717180972
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 1717180972
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_43
timestamp 1717180972
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1717180972
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1717180972
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1717180972
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1717180972
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_97
timestamp 1717180972
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_101
timestamp 1717180972
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1717180972
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1717180972
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1717180972
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1717180972
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_43
timestamp 1717180972
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_55
timestamp 1717180972
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1717180972
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1717180972
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_29
timestamp 1717180972
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1717180972
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1717180972
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_77
timestamp 1717180972
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_96
timestamp 1717180972
transform 1 0 9936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1717180972
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 1717180972
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_40
timestamp 1717180972
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_44
timestamp 1717180972
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_68
timestamp 1717180972
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_76
timestamp 1717180972
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1717180972
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1717180972
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_99
timestamp 1717180972
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1717180972
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1717180972
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 1717180972
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1717180972
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1717180972
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_61
timestamp 1717180972
transform 1 0 6716 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_69
timestamp 1717180972
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_75
timestamp 1717180972
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1717180972
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1717180972
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1717180972
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1717180972
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_32
timestamp 1717180972
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_66
timestamp 1717180972
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1717180972
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1717180972
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_26
timestamp 1717180972
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_49
timestamp 1717180972
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 1717180972
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_86
timestamp 1717180972
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_101
timestamp 1717180972
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1717180972
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_12
timestamp 1717180972
transform 1 0 2208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_20
timestamp 1717180972
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1717180972
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 1717180972
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1717180972
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1717180972
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_100
timestamp 1717180972
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1717180972
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_25
timestamp 1717180972
transform 1 0 3404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_29
timestamp 1717180972
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1717180972
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1717180972
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1717180972
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_62
timestamp 1717180972
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_71
timestamp 1717180972
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_90
timestamp 1717180972
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1717180972
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1717180972
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1717180972
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1717180972
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1717180972
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_42
timestamp 1717180972
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_52
timestamp 1717180972
transform 1 0 5888 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_58
timestamp 1717180972
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_70
timestamp 1717180972
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1717180972
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1717180972
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1717180972
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1717180972
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_44
timestamp 1717180972
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1717180972
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_72
timestamp 1717180972
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_82
timestamp 1717180972
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1717180972
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1717180972
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1717180972
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1717180972
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1717180972
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_96
timestamp 1717180972
transform 1 0 9936 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_6
timestamp 1717180972
transform 1 0 1656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_12
timestamp 1717180972
transform 1 0 2208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_28
timestamp 1717180972
transform 1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1717180972
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_71
timestamp 1717180972
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_87
timestamp 1717180972
transform 1 0 9108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1717180972
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_15
timestamp 1717180972
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1717180972
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_29
timestamp 1717180972
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_40
timestamp 1717180972
transform 1 0 4784 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_52
timestamp 1717180972
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_57
timestamp 1717180972
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_68
timestamp 1717180972
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1717180972
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1717180972
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_92
timestamp 1717180972
transform 1 0 9568 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_100
timestamp 1717180972
transform 1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1717180972
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1717180972
transform -1 0 8740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1717180972
transform 1 0 7268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1717180972
transform -1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1717180972
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1717180972
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1717180972
transform -1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1717180972
transform -1 0 4784 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1717180972
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1717180972
transform -1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1717180972
transform -1 0 9936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1717180972
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1717180972
transform -1 0 3128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1717180972
transform -1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold17
timestamp 1717180972
transform -1 0 5336 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1717180972
transform 1 0 4048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  hold20
timestamp 1717180972
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1717180972
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold22
timestamp 1717180972
transform 1 0 4140 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1717180972
transform 1 0 5152 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1717180972
transform -1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold25
timestamp 1717180972
transform -1 0 4140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1717180972
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1717180972
transform -1 0 10396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1717180972
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1717180972
transform -1 0 8648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1717180972
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1717180972
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1717180972
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1717180972
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1717180972
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1717180972
transform 1 0 9016 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1717180972
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1717180972
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1717180972
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1717180972
transform -1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1717180972
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1717180972
transform -1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1717180972
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1717180972
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1717180972
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1717180972
transform -1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1717180972
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1717180972
transform -1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1717180972
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1717180972
transform -1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1717180972
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1717180972
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1717180972
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1717180972
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1717180972
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1717180972
transform -1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1717180972
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1717180972
transform -1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1717180972
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1717180972
transform -1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1717180972
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1717180972
transform -1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1717180972
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1717180972
transform -1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1717180972
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1717180972
transform -1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1717180972
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1717180972
transform -1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1717180972
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1717180972
transform -1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717180972
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1717180972
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1717180972
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1717180972
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1717180972
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1717180972
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1717180972
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1717180972
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1717180972
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1717180972
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1717180972
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1717180972
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1717180972
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1717180972
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1717180972
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1717180972
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1717180972
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1717180972
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1717180972
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1717180972
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1717180972
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1717180972
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1717180972
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1717180972
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1717180972
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1717180972
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1717180972
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1717180972
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 3358 2128 3678 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5773 2128 6093 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8188 2128 8508 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10603 2128 10923 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2151 2128 2471 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4566 2128 4886 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6981 2128 7301 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9396 2128 9716 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 11154 3272 11954 3392 0 FreeSans 480 0 0 0 percentage[0]
port 3 nsew signal input
flabel metal3 s 11154 10344 11954 10464 0 FreeSans 480 0 0 0 percentage[1]
port 4 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 s_in_lines[0]
port 5 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 s_in_lines[1]
port 6 nsew signal input
flabel metal2 s 2962 13298 3018 14098 0 FreeSans 224 90 0 0 s_out_lines[0]
port 7 nsew signal tristate
flabel metal2 s 8942 13298 8998 14098 0 FreeSans 224 90 0 0 s_out_lines[1]
port 8 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 start
port 9 nsew signal input
rlabel via1 6013 10880 6013 10880 0 VGND
rlabel metal1 5934 11424 5934 11424 0 VPWR
rlabel metal2 7774 7684 7774 7684 0 CTRLPTH1.done
rlabel metal1 7590 8602 7590 8602 0 CTRLPTH1.state\[0\]
rlabel metal1 5428 8942 5428 8942 0 CTRLPTH1.state\[1\]
rlabel metal1 7360 10574 7360 10574 0 CTRLPTH1.state\[2\]
rlabel metal1 10626 9010 10626 9010 0 DTPTH1.PS1.count\[0\]
rlabel metal2 9338 8058 9338 8058 0 DTPTH1.PS1.count\[1\]
rlabel metal1 3818 6732 3818 6732 0 DTPTH1.RS1.RNG1.TFF1.Q
rlabel metal1 4048 8466 4048 8466 0 DTPTH1.RS1.RNG1.TFF2.Q
rlabel metal1 5428 6834 5428 6834 0 DTPTH1.RS1.RNG1.TFF3.Q
rlabel metal2 4002 5508 4002 5508 0 DTPTH1.RS1.RNG1.TFF4.Q
rlabel metal1 3956 4658 3956 4658 0 DTPTH1.RS1.RNG1.TFF5.Q
rlabel metal1 5198 3434 5198 3434 0 DTPTH1.RS1.RNG1.TFF6.Q
rlabel metal1 4370 3468 4370 3468 0 DTPTH1.RS1.RNG1.TFF7.Q
rlabel metal1 4738 6154 4738 6154 0 DTPTH1.RS1.RNG1.b0
rlabel metal1 6118 5270 6118 5270 0 DTPTH1.RS1.RNG1.b1
rlabel metal1 5106 4046 5106 4046 0 DTPTH1.RS1.RNG1.b2
rlabel metal1 7866 4114 7866 4114 0 DTPTH1.RS1.RNG1.r_num\[0\]
rlabel metal1 8786 3434 8786 3434 0 DTPTH1.RS1.RNG1.r_num\[1\]
rlabel metal1 7866 5882 7866 5882 0 DTPTH1.RS1.RNG1.r_num\[2\]
rlabel metal1 10212 7378 10212 7378 0 DTPTH1.RS1.counter\[0\]
rlabel metal1 9522 6868 9522 6868 0 DTPTH1.RS1.counter\[1\]
rlabel metal1 10120 4658 10120 4658 0 DTPTH1.RS1.s_comb\[0\]
rlabel metal1 10212 3706 10212 3706 0 DTPTH1.RS1.s_comb\[1\]
rlabel metal2 8694 4182 8694 4182 0 DTPTH1.RS1.s_comb\[2\]
rlabel metal1 9292 2482 9292 2482 0 DTPTH1.RS1.s_comb\[3\]
rlabel metal1 5435 7378 5435 7378 0 _000_
rlabel metal1 4646 9486 4646 9486 0 _001_
rlabel metal1 2944 3026 2944 3026 0 _002_
rlabel metal1 6568 7378 6568 7378 0 _003_
rlabel metal1 9752 4794 9752 4794 0 _004_
rlabel metal1 9246 3060 9246 3060 0 _005_
rlabel metal1 7268 4250 7268 4250 0 _006_
rlabel metal1 8004 2618 8004 2618 0 _007_
rlabel metal1 4048 2346 4048 2346 0 _008_
rlabel metal1 2484 5134 2484 5134 0 _009_
rlabel metal1 3864 5746 3864 5746 0 _010_
rlabel metal1 3036 7922 3036 7922 0 _011_
rlabel metal1 1748 8058 1748 8058 0 _012_
rlabel metal2 1978 7140 1978 7140 0 _013_
rlabel metal1 8970 6392 8970 6392 0 _014_
rlabel metal2 7774 6562 7774 6562 0 _015_
rlabel metal1 3986 9962 3986 9962 0 _016_
rlabel metal1 5581 10710 5581 10710 0 _017_
rlabel metal2 6578 9826 6578 9826 0 _018_
rlabel metal1 9425 9622 9425 9622 0 _019_
rlabel metal1 8178 8466 8178 8466 0 _020_
rlabel metal1 6990 9554 6990 9554 0 _021_
rlabel metal1 3956 9010 3956 9010 0 _022_
rlabel metal1 7130 10642 7130 10642 0 _023_
rlabel metal1 9890 10064 9890 10064 0 _024_
rlabel metal1 8372 9554 8372 9554 0 _025_
rlabel metal2 7406 10302 7406 10302 0 _026_
rlabel metal1 7912 8874 7912 8874 0 _027_
rlabel metal2 9982 6426 9982 6426 0 _028_
rlabel metal1 7544 7174 7544 7174 0 _029_
rlabel metal1 5934 7412 5934 7412 0 _030_
rlabel metal1 9062 4250 9062 4250 0 _031_
rlabel metal1 8970 8874 8970 8874 0 _032_
rlabel metal1 7958 2550 7958 2550 0 _033_
rlabel metal1 7222 3094 7222 3094 0 _034_
rlabel metal1 8188 2414 8188 2414 0 _035_
rlabel metal1 2346 5746 2346 5746 0 _036_
rlabel metal2 1886 6358 1886 6358 0 _037_
rlabel metal1 7958 7310 7958 7310 0 _038_
rlabel metal1 9384 7514 9384 7514 0 _039_
rlabel metal1 10074 6834 10074 6834 0 _040_
rlabel metal2 10166 6698 10166 6698 0 _041_
rlabel metal1 9936 5882 9936 5882 0 _042_
rlabel metal1 8648 7446 8648 7446 0 _043_
rlabel metal1 8648 7514 8648 7514 0 _044_
rlabel metal1 5750 10608 5750 10608 0 _045_
rlabel metal1 3542 10234 3542 10234 0 _046_
rlabel metal2 8418 10472 8418 10472 0 _047_
rlabel metal2 8142 10472 8142 10472 0 _048_
rlabel metal3 1671 3332 1671 3332 0 clk
rlabel metal1 6440 6630 6440 6630 0 clknet_0_clk
rlabel metal1 1794 3570 1794 3570 0 clknet_1_0__leaf_clk
rlabel metal1 1702 7446 1702 7446 0 clknet_1_1__leaf_clk
rlabel metal1 9936 10234 9936 10234 0 net1
rlabel metal1 7498 4080 7498 4080 0 net10
rlabel metal1 7677 3434 7677 3434 0 net11
rlabel metal1 8740 2414 8740 2414 0 net12
rlabel metal2 5566 9690 5566 9690 0 net13
rlabel metal2 6026 9146 6026 9146 0 net14
rlabel metal1 4363 2346 4363 2346 0 net15
rlabel metal1 4738 9554 4738 9554 0 net16
rlabel metal2 3266 10608 3266 10608 0 net17
rlabel metal1 5014 9146 5014 9146 0 net18
rlabel metal1 9614 4590 9614 4590 0 net19
rlabel metal1 9200 10030 9200 10030 0 net2
rlabel metal1 9011 5270 9011 5270 0 net20
rlabel metal1 3680 3026 3680 3026 0 net21
rlabel metal1 2162 3162 2162 3162 0 net22
rlabel metal1 7360 9486 7360 9486 0 net23
rlabel metal1 3312 5746 3312 5746 0 net24
rlabel metal1 5474 5304 5474 5304 0 net25
rlabel metal2 5290 4760 5290 4760 0 net26
rlabel metal1 3450 6970 3450 6970 0 net27
rlabel metal2 5842 5916 5842 5916 0 net28
rlabel metal1 3818 4114 3818 4114 0 net29
rlabel metal1 2990 2618 2990 2618 0 net3
rlabel metal1 5651 3706 5651 3706 0 net30
rlabel metal1 3956 3706 3956 3706 0 net31
rlabel metal1 3726 7922 3726 7922 0 net32
rlabel metal1 9752 8942 9752 8942 0 net33
rlabel metal1 8510 6290 8510 6290 0 net34
rlabel metal1 8786 6970 8786 6970 0 net35
rlabel metal1 7958 6358 7958 6358 0 net36
rlabel metal1 8464 2278 8464 2278 0 net4
rlabel metal1 1610 10132 1610 10132 0 net5
rlabel metal2 3174 10914 3174 10914 0 net6
rlabel metal1 9108 10778 9108 10778 0 net7
rlabel metal1 8464 2822 8464 2822 0 net8
rlabel metal2 9890 3298 9890 3298 0 net9
rlabel metal1 10672 3026 10672 3026 0 percentage[0]
rlabel metal1 10672 10642 10672 10642 0 percentage[1]
rlabel metal2 2990 1588 2990 1588 0 s_in_lines[0]
rlabel metal2 8970 1027 8970 1027 0 s_in_lines[1]
rlabel metal1 3128 11322 3128 11322 0 s_out_lines[0]
rlabel metal1 9108 11322 9108 11322 0 s_out_lines[1]
rlabel metal3 820 10404 820 10404 0 start
<< properties >>
string FIXED_BBOX 0 0 11954 14098
<< end >>
